magic
tech sky130A
magscale 1 2
timestamp 1693602505
<< nwell >>
rect 1066 349509 558846 349830
rect 1066 348421 558846 348987
rect 1066 347333 558846 347899
rect 1066 346245 558846 346811
rect 1066 345157 558846 345723
rect 1066 344069 558846 344635
rect 1066 342981 558846 343547
rect 1066 341893 558846 342459
rect 1066 340805 558846 341371
rect 1066 339717 558846 340283
rect 1066 338629 558846 339195
rect 1066 337541 558846 338107
rect 1066 336453 558846 337019
rect 1066 335365 558846 335931
rect 1066 334277 558846 334843
rect 1066 333189 558846 333755
rect 1066 332101 558846 332667
rect 1066 331013 558846 331579
rect 1066 329925 558846 330491
rect 1066 328837 558846 329403
rect 1066 327749 558846 328315
rect 1066 326661 558846 327227
rect 1066 325573 558846 326139
rect 1066 324485 558846 325051
rect 1066 323397 558846 323963
rect 1066 322309 558846 322875
rect 1066 321221 558846 321787
rect 1066 320133 558846 320699
rect 1066 319045 558846 319611
rect 1066 317957 558846 318523
rect 1066 316869 558846 317435
rect 1066 315781 558846 316347
rect 1066 314693 558846 315259
rect 1066 313605 558846 314171
rect 1066 312517 558846 313083
rect 1066 311429 558846 311995
rect 1066 310341 558846 310907
rect 1066 309253 558846 309819
rect 1066 308165 558846 308731
rect 1066 307077 558846 307643
rect 1066 305989 558846 306555
rect 1066 304901 558846 305467
rect 1066 303813 558846 304379
rect 1066 302725 558846 303291
rect 1066 301637 558846 302203
rect 1066 300549 558846 301115
rect 1066 299461 558846 300027
rect 1066 298373 558846 298939
rect 1066 297285 558846 297851
rect 1066 296197 558846 296763
rect 1066 295109 558846 295675
rect 1066 294021 558846 294587
rect 1066 292933 558846 293499
rect 1066 291845 558846 292411
rect 1066 290757 558846 291323
rect 1066 289669 558846 290235
rect 1066 288581 558846 289147
rect 1066 287493 558846 288059
rect 1066 286405 558846 286971
rect 1066 285317 558846 285883
rect 1066 284229 558846 284795
rect 1066 283141 558846 283707
rect 1066 282053 558846 282619
rect 1066 280965 558846 281531
rect 1066 279877 558846 280443
rect 1066 278789 558846 279355
rect 1066 277701 558846 278267
rect 1066 276613 558846 277179
rect 1066 275525 558846 276091
rect 1066 274437 558846 275003
rect 1066 273349 558846 273915
rect 1066 272261 558846 272827
rect 1066 271173 558846 271739
rect 1066 270085 558846 270651
rect 1066 268997 558846 269563
rect 1066 267909 558846 268475
rect 1066 266821 558846 267387
rect 1066 265733 558846 266299
rect 1066 264645 558846 265211
rect 1066 263557 558846 264123
rect 1066 262469 558846 263035
rect 1066 261381 558846 261947
rect 1066 260293 558846 260859
rect 1066 259205 558846 259771
rect 1066 258117 558846 258683
rect 1066 257029 558846 257595
rect 1066 255941 558846 256507
rect 1066 254853 558846 255419
rect 1066 253765 558846 254331
rect 1066 252677 558846 253243
rect 1066 251589 558846 252155
rect 1066 250501 558846 251067
rect 1066 249413 558846 249979
rect 1066 248325 558846 248891
rect 1066 247237 558846 247803
rect 1066 246149 558846 246715
rect 1066 245061 558846 245627
rect 1066 243973 558846 244539
rect 1066 242885 558846 243451
rect 1066 241797 558846 242363
rect 1066 240709 558846 241275
rect 1066 239621 558846 240187
rect 1066 238533 558846 239099
rect 1066 237445 558846 238011
rect 1066 236357 558846 236923
rect 1066 235269 558846 235835
rect 1066 234181 558846 234747
rect 1066 233093 558846 233659
rect 1066 232005 558846 232571
rect 1066 230917 558846 231483
rect 1066 229829 558846 230395
rect 1066 228741 558846 229307
rect 1066 227653 558846 228219
rect 1066 226565 558846 227131
rect 1066 225477 558846 226043
rect 1066 224389 558846 224955
rect 1066 223301 558846 223867
rect 1066 222213 558846 222779
rect 1066 221125 558846 221691
rect 1066 220037 558846 220603
rect 1066 218949 558846 219515
rect 1066 217861 558846 218427
rect 1066 216773 558846 217339
rect 1066 215685 558846 216251
rect 1066 214597 558846 215163
rect 1066 213509 558846 214075
rect 1066 212421 558846 212987
rect 1066 211333 558846 211899
rect 1066 210245 558846 210811
rect 1066 209157 558846 209723
rect 1066 208069 558846 208635
rect 1066 206981 558846 207547
rect 1066 205893 558846 206459
rect 1066 204805 558846 205371
rect 1066 203717 558846 204283
rect 1066 202629 558846 203195
rect 1066 201541 558846 202107
rect 1066 200453 558846 201019
rect 1066 199365 558846 199931
rect 1066 198277 558846 198843
rect 1066 197189 558846 197755
rect 1066 196101 558846 196667
rect 1066 195013 558846 195579
rect 1066 193925 558846 194491
rect 1066 192837 558846 193403
rect 1066 191749 558846 192315
rect 1066 190661 558846 191227
rect 1066 189573 558846 190139
rect 1066 188485 558846 189051
rect 1066 187397 558846 187963
rect 1066 186309 558846 186875
rect 1066 185221 558846 185787
rect 1066 184133 558846 184699
rect 1066 183045 558846 183611
rect 1066 181957 558846 182523
rect 1066 180869 558846 181435
rect 1066 179781 558846 180347
rect 1066 178693 558846 179259
rect 1066 177605 558846 178171
rect 1066 176517 558846 177083
rect 1066 175429 558846 175995
rect 1066 174341 558846 174907
rect 1066 173253 558846 173819
rect 1066 172165 558846 172731
rect 1066 171077 558846 171643
rect 1066 169989 558846 170555
rect 1066 168901 558846 169467
rect 1066 167813 558846 168379
rect 1066 166725 558846 167291
rect 1066 165637 558846 166203
rect 1066 164549 558846 165115
rect 1066 163461 558846 164027
rect 1066 162373 558846 162939
rect 1066 161285 558846 161851
rect 1066 160197 558846 160763
rect 1066 159109 558846 159675
rect 1066 158021 558846 158587
rect 1066 156933 558846 157499
rect 1066 155845 558846 156411
rect 1066 154757 558846 155323
rect 1066 153669 558846 154235
rect 1066 152581 558846 153147
rect 1066 151493 558846 152059
rect 1066 150405 558846 150971
rect 1066 149317 558846 149883
rect 1066 148229 558846 148795
rect 1066 147141 558846 147707
rect 1066 146053 558846 146619
rect 1066 144965 558846 145531
rect 1066 143877 558846 144443
rect 1066 142789 558846 143355
rect 1066 141701 558846 142267
rect 1066 140613 558846 141179
rect 1066 139525 558846 140091
rect 1066 138437 558846 139003
rect 1066 137349 558846 137915
rect 1066 136261 558846 136827
rect 1066 135173 558846 135739
rect 1066 134085 558846 134651
rect 1066 132997 558846 133563
rect 1066 131909 558846 132475
rect 1066 130821 558846 131387
rect 1066 129733 558846 130299
rect 1066 128645 558846 129211
rect 1066 127557 558846 128123
rect 1066 126469 558846 127035
rect 1066 125381 558846 125947
rect 1066 124293 558846 124859
rect 1066 123205 558846 123771
rect 1066 122117 558846 122683
rect 1066 121029 558846 121595
rect 1066 119941 558846 120507
rect 1066 118853 558846 119419
rect 1066 117765 558846 118331
rect 1066 116677 558846 117243
rect 1066 115589 558846 116155
rect 1066 114501 558846 115067
rect 1066 113413 558846 113979
rect 1066 112325 558846 112891
rect 1066 111237 558846 111803
rect 1066 110149 558846 110715
rect 1066 109061 558846 109627
rect 1066 107973 558846 108539
rect 1066 106885 558846 107451
rect 1066 105797 558846 106363
rect 1066 104709 558846 105275
rect 1066 103621 558846 104187
rect 1066 102533 558846 103099
rect 1066 101445 558846 102011
rect 1066 100357 558846 100923
rect 1066 99269 558846 99835
rect 1066 98181 558846 98747
rect 1066 97093 558846 97659
rect 1066 96005 558846 96571
rect 1066 94917 558846 95483
rect 1066 93829 558846 94395
rect 1066 92741 558846 93307
rect 1066 91653 558846 92219
rect 1066 90565 558846 91131
rect 1066 89477 558846 90043
rect 1066 88389 558846 88955
rect 1066 87301 558846 87867
rect 1066 86213 558846 86779
rect 1066 85125 558846 85691
rect 1066 84037 558846 84603
rect 1066 82949 558846 83515
rect 1066 81861 558846 82427
rect 1066 80773 558846 81339
rect 1066 79685 558846 80251
rect 1066 78597 558846 79163
rect 1066 77509 558846 78075
rect 1066 76421 558846 76987
rect 1066 75333 558846 75899
rect 1066 74245 558846 74811
rect 1066 73157 558846 73723
rect 1066 72069 558846 72635
rect 1066 70981 558846 71547
rect 1066 69893 558846 70459
rect 1066 68805 558846 69371
rect 1066 67717 558846 68283
rect 1066 66629 558846 67195
rect 1066 65541 558846 66107
rect 1066 64453 558846 65019
rect 1066 63365 558846 63931
rect 1066 62277 558846 62843
rect 1066 61189 558846 61755
rect 1066 60101 558846 60667
rect 1066 59013 558846 59579
rect 1066 57925 558846 58491
rect 1066 56837 558846 57403
rect 1066 55749 558846 56315
rect 1066 54661 558846 55227
rect 1066 53573 558846 54139
rect 1066 52485 558846 53051
rect 1066 51397 558846 51963
rect 1066 50309 558846 50875
rect 1066 49221 558846 49787
rect 1066 48133 558846 48699
rect 1066 47045 558846 47611
rect 1066 45957 558846 46523
rect 1066 44869 558846 45435
rect 1066 43781 558846 44347
rect 1066 42693 558846 43259
rect 1066 41605 558846 42171
rect 1066 40517 558846 41083
rect 1066 39429 558846 39995
rect 1066 38341 558846 38907
rect 1066 37253 558846 37819
rect 1066 36165 558846 36731
rect 1066 35077 558846 35643
rect 1066 33989 558846 34555
rect 1066 32901 558846 33467
rect 1066 31813 558846 32379
rect 1066 30725 558846 31291
rect 1066 29637 558846 30203
rect 1066 28549 558846 29115
rect 1066 27461 558846 28027
rect 1066 26373 558846 26939
rect 1066 25285 558846 25851
rect 1066 24197 558846 24763
rect 1066 23109 558846 23675
rect 1066 22021 558846 22587
rect 1066 20933 558846 21499
rect 1066 19845 558846 20411
rect 1066 18757 558846 19323
rect 1066 17669 558846 18235
rect 1066 16581 558846 17147
rect 1066 15493 558846 16059
rect 1066 14405 558846 14971
rect 1066 13317 558846 13883
rect 1066 12229 558846 12795
rect 1066 11141 558846 11707
rect 1066 10053 558846 10619
rect 1066 8965 558846 9531
rect 1066 7877 558846 8443
rect 1066 6789 558846 7355
rect 1066 5701 558846 6267
rect 1066 4613 558846 5179
rect 1066 3525 558846 4091
rect 1066 2437 558846 3003
<< obsli1 >>
rect 1104 2159 558808 349809
<< obsm1 >>
rect 1104 144 558808 349840
<< metal2 >>
rect 7010 0 7066 800
rect 11242 0 11298 800
rect 15474 0 15530 800
rect 19706 0 19762 800
rect 23938 0 23994 800
rect 28170 0 28226 800
rect 32402 0 32458 800
rect 36634 0 36690 800
rect 40866 0 40922 800
rect 45098 0 45154 800
rect 49330 0 49386 800
rect 53562 0 53618 800
rect 57794 0 57850 800
rect 62026 0 62082 800
rect 66258 0 66314 800
rect 70490 0 70546 800
rect 74722 0 74778 800
rect 78954 0 79010 800
rect 83186 0 83242 800
rect 87418 0 87474 800
rect 91650 0 91706 800
rect 95882 0 95938 800
rect 100114 0 100170 800
rect 104346 0 104402 800
rect 108578 0 108634 800
rect 112810 0 112866 800
rect 117042 0 117098 800
rect 121274 0 121330 800
rect 125506 0 125562 800
rect 129738 0 129794 800
rect 133970 0 134026 800
rect 138202 0 138258 800
rect 142434 0 142490 800
rect 146666 0 146722 800
rect 150898 0 150954 800
rect 155130 0 155186 800
rect 159362 0 159418 800
rect 163594 0 163650 800
rect 167826 0 167882 800
rect 172058 0 172114 800
rect 176290 0 176346 800
rect 180522 0 180578 800
rect 184754 0 184810 800
rect 188986 0 189042 800
rect 193218 0 193274 800
rect 197450 0 197506 800
rect 201682 0 201738 800
rect 205914 0 205970 800
rect 210146 0 210202 800
rect 214378 0 214434 800
rect 218610 0 218666 800
rect 222842 0 222898 800
rect 227074 0 227130 800
rect 231306 0 231362 800
rect 235538 0 235594 800
rect 239770 0 239826 800
rect 244002 0 244058 800
rect 248234 0 248290 800
rect 252466 0 252522 800
rect 256698 0 256754 800
rect 260930 0 260986 800
rect 265162 0 265218 800
rect 269394 0 269450 800
rect 273626 0 273682 800
rect 277858 0 277914 800
rect 282090 0 282146 800
rect 286322 0 286378 800
rect 290554 0 290610 800
rect 294786 0 294842 800
rect 299018 0 299074 800
rect 303250 0 303306 800
rect 307482 0 307538 800
rect 311714 0 311770 800
rect 315946 0 316002 800
rect 320178 0 320234 800
rect 324410 0 324466 800
rect 328642 0 328698 800
rect 332874 0 332930 800
rect 337106 0 337162 800
rect 341338 0 341394 800
rect 345570 0 345626 800
rect 349802 0 349858 800
rect 354034 0 354090 800
rect 358266 0 358322 800
rect 362498 0 362554 800
rect 366730 0 366786 800
rect 370962 0 371018 800
rect 375194 0 375250 800
rect 379426 0 379482 800
rect 383658 0 383714 800
rect 387890 0 387946 800
rect 392122 0 392178 800
rect 396354 0 396410 800
rect 400586 0 400642 800
rect 404818 0 404874 800
rect 409050 0 409106 800
rect 413282 0 413338 800
rect 417514 0 417570 800
rect 421746 0 421802 800
rect 425978 0 426034 800
rect 430210 0 430266 800
rect 434442 0 434498 800
rect 438674 0 438730 800
rect 442906 0 442962 800
rect 447138 0 447194 800
rect 451370 0 451426 800
rect 455602 0 455658 800
rect 459834 0 459890 800
rect 464066 0 464122 800
rect 468298 0 468354 800
rect 472530 0 472586 800
rect 476762 0 476818 800
rect 480994 0 481050 800
rect 485226 0 485282 800
rect 489458 0 489514 800
rect 493690 0 493746 800
rect 497922 0 497978 800
rect 502154 0 502210 800
rect 506386 0 506442 800
rect 510618 0 510674 800
rect 514850 0 514906 800
rect 519082 0 519138 800
rect 523314 0 523370 800
rect 527546 0 527602 800
rect 531778 0 531834 800
rect 536010 0 536066 800
rect 540242 0 540298 800
rect 544474 0 544530 800
rect 548706 0 548762 800
rect 552938 0 552994 800
<< obsm2 >>
rect 4214 856 557482 349829
rect 4214 31 6954 856
rect 7122 31 11186 856
rect 11354 31 15418 856
rect 15586 31 19650 856
rect 19818 31 23882 856
rect 24050 31 28114 856
rect 28282 31 32346 856
rect 32514 31 36578 856
rect 36746 31 40810 856
rect 40978 31 45042 856
rect 45210 31 49274 856
rect 49442 31 53506 856
rect 53674 31 57738 856
rect 57906 31 61970 856
rect 62138 31 66202 856
rect 66370 31 70434 856
rect 70602 31 74666 856
rect 74834 31 78898 856
rect 79066 31 83130 856
rect 83298 31 87362 856
rect 87530 31 91594 856
rect 91762 31 95826 856
rect 95994 31 100058 856
rect 100226 31 104290 856
rect 104458 31 108522 856
rect 108690 31 112754 856
rect 112922 31 116986 856
rect 117154 31 121218 856
rect 121386 31 125450 856
rect 125618 31 129682 856
rect 129850 31 133914 856
rect 134082 31 138146 856
rect 138314 31 142378 856
rect 142546 31 146610 856
rect 146778 31 150842 856
rect 151010 31 155074 856
rect 155242 31 159306 856
rect 159474 31 163538 856
rect 163706 31 167770 856
rect 167938 31 172002 856
rect 172170 31 176234 856
rect 176402 31 180466 856
rect 180634 31 184698 856
rect 184866 31 188930 856
rect 189098 31 193162 856
rect 193330 31 197394 856
rect 197562 31 201626 856
rect 201794 31 205858 856
rect 206026 31 210090 856
rect 210258 31 214322 856
rect 214490 31 218554 856
rect 218722 31 222786 856
rect 222954 31 227018 856
rect 227186 31 231250 856
rect 231418 31 235482 856
rect 235650 31 239714 856
rect 239882 31 243946 856
rect 244114 31 248178 856
rect 248346 31 252410 856
rect 252578 31 256642 856
rect 256810 31 260874 856
rect 261042 31 265106 856
rect 265274 31 269338 856
rect 269506 31 273570 856
rect 273738 31 277802 856
rect 277970 31 282034 856
rect 282202 31 286266 856
rect 286434 31 290498 856
rect 290666 31 294730 856
rect 294898 31 298962 856
rect 299130 31 303194 856
rect 303362 31 307426 856
rect 307594 31 311658 856
rect 311826 31 315890 856
rect 316058 31 320122 856
rect 320290 31 324354 856
rect 324522 31 328586 856
rect 328754 31 332818 856
rect 332986 31 337050 856
rect 337218 31 341282 856
rect 341450 31 345514 856
rect 345682 31 349746 856
rect 349914 31 353978 856
rect 354146 31 358210 856
rect 358378 31 362442 856
rect 362610 31 366674 856
rect 366842 31 370906 856
rect 371074 31 375138 856
rect 375306 31 379370 856
rect 379538 31 383602 856
rect 383770 31 387834 856
rect 388002 31 392066 856
rect 392234 31 396298 856
rect 396466 31 400530 856
rect 400698 31 404762 856
rect 404930 31 408994 856
rect 409162 31 413226 856
rect 413394 31 417458 856
rect 417626 31 421690 856
rect 421858 31 425922 856
rect 426090 31 430154 856
rect 430322 31 434386 856
rect 434554 31 438618 856
rect 438786 31 442850 856
rect 443018 31 447082 856
rect 447250 31 451314 856
rect 451482 31 455546 856
rect 455714 31 459778 856
rect 459946 31 464010 856
rect 464178 31 468242 856
rect 468410 31 472474 856
rect 472642 31 476706 856
rect 476874 31 480938 856
rect 481106 31 485170 856
rect 485338 31 489402 856
rect 489570 31 493634 856
rect 493802 31 497866 856
rect 498034 31 502098 856
rect 502266 31 506330 856
rect 506498 31 510562 856
rect 510730 31 514794 856
rect 514962 31 519026 856
rect 519194 31 523258 856
rect 523426 31 527490 856
rect 527658 31 531722 856
rect 531890 31 535954 856
rect 536122 31 540186 856
rect 540354 31 544418 856
rect 544586 31 548650 856
rect 548818 31 552882 856
rect 553050 31 557482 856
<< obsm3 >>
rect 4210 35 557486 349825
<< metal4 >>
rect 4208 2128 4528 349840
rect 19568 2128 19888 349840
rect 34928 2128 35248 349840
rect 50288 2128 50608 349840
rect 65648 2128 65968 349840
rect 81008 2128 81328 349840
rect 96368 2128 96688 349840
rect 111728 2128 112048 349840
rect 127088 2128 127408 349840
rect 142448 2128 142768 349840
rect 157808 2128 158128 349840
rect 173168 2128 173488 349840
rect 188528 2128 188848 349840
rect 203888 2128 204208 349840
rect 219248 2128 219568 349840
rect 234608 2128 234928 349840
rect 249968 2128 250288 349840
rect 265328 2128 265648 349840
rect 280688 2128 281008 349840
rect 296048 2128 296368 349840
rect 311408 2128 311728 349840
rect 326768 2128 327088 349840
rect 342128 2128 342448 349840
rect 357488 2128 357808 349840
rect 372848 2128 373168 349840
rect 388208 2128 388528 349840
rect 403568 2128 403888 349840
rect 418928 2128 419248 349840
rect 434288 2128 434608 349840
rect 449648 2128 449968 349840
rect 465008 2128 465328 349840
rect 480368 2128 480688 349840
rect 495728 2128 496048 349840
rect 511088 2128 511408 349840
rect 526448 2128 526768 349840
rect 541808 2128 542128 349840
rect 557168 2128 557488 349840
<< obsm4 >>
rect 191603 2048 203808 29613
rect 204288 2048 219168 29613
rect 219648 2048 234528 29613
rect 235008 2048 249888 29613
rect 250368 2048 265248 29613
rect 265728 2048 278149 29613
rect 191603 35 278149 2048
<< labels >>
rlabel metal2 s 11242 0 11298 800 6 la_data_in[0]
port 1 nsew signal input
rlabel metal2 s 95882 0 95938 800 6 la_data_in[10]
port 2 nsew signal input
rlabel metal2 s 104346 0 104402 800 6 la_data_in[11]
port 3 nsew signal input
rlabel metal2 s 112810 0 112866 800 6 la_data_in[12]
port 4 nsew signal input
rlabel metal2 s 121274 0 121330 800 6 la_data_in[13]
port 5 nsew signal input
rlabel metal2 s 129738 0 129794 800 6 la_data_in[14]
port 6 nsew signal input
rlabel metal2 s 138202 0 138258 800 6 la_data_in[15]
port 7 nsew signal input
rlabel metal2 s 146666 0 146722 800 6 la_data_in[16]
port 8 nsew signal input
rlabel metal2 s 155130 0 155186 800 6 la_data_in[17]
port 9 nsew signal input
rlabel metal2 s 163594 0 163650 800 6 la_data_in[18]
port 10 nsew signal input
rlabel metal2 s 172058 0 172114 800 6 la_data_in[19]
port 11 nsew signal input
rlabel metal2 s 19706 0 19762 800 6 la_data_in[1]
port 12 nsew signal input
rlabel metal2 s 180522 0 180578 800 6 la_data_in[20]
port 13 nsew signal input
rlabel metal2 s 188986 0 189042 800 6 la_data_in[21]
port 14 nsew signal input
rlabel metal2 s 197450 0 197506 800 6 la_data_in[22]
port 15 nsew signal input
rlabel metal2 s 205914 0 205970 800 6 la_data_in[23]
port 16 nsew signal input
rlabel metal2 s 214378 0 214434 800 6 la_data_in[24]
port 17 nsew signal input
rlabel metal2 s 222842 0 222898 800 6 la_data_in[25]
port 18 nsew signal input
rlabel metal2 s 231306 0 231362 800 6 la_data_in[26]
port 19 nsew signal input
rlabel metal2 s 239770 0 239826 800 6 la_data_in[27]
port 20 nsew signal input
rlabel metal2 s 248234 0 248290 800 6 la_data_in[28]
port 21 nsew signal input
rlabel metal2 s 256698 0 256754 800 6 la_data_in[29]
port 22 nsew signal input
rlabel metal2 s 28170 0 28226 800 6 la_data_in[2]
port 23 nsew signal input
rlabel metal2 s 265162 0 265218 800 6 la_data_in[30]
port 24 nsew signal input
rlabel metal2 s 273626 0 273682 800 6 la_data_in[31]
port 25 nsew signal input
rlabel metal2 s 282090 0 282146 800 6 la_data_in[32]
port 26 nsew signal input
rlabel metal2 s 290554 0 290610 800 6 la_data_in[33]
port 27 nsew signal input
rlabel metal2 s 294786 0 294842 800 6 la_data_in[34]
port 28 nsew signal input
rlabel metal2 s 299018 0 299074 800 6 la_data_in[35]
port 29 nsew signal input
rlabel metal2 s 303250 0 303306 800 6 la_data_in[36]
port 30 nsew signal input
rlabel metal2 s 307482 0 307538 800 6 la_data_in[37]
port 31 nsew signal input
rlabel metal2 s 311714 0 311770 800 6 la_data_in[38]
port 32 nsew signal input
rlabel metal2 s 315946 0 316002 800 6 la_data_in[39]
port 33 nsew signal input
rlabel metal2 s 36634 0 36690 800 6 la_data_in[3]
port 34 nsew signal input
rlabel metal2 s 320178 0 320234 800 6 la_data_in[40]
port 35 nsew signal input
rlabel metal2 s 324410 0 324466 800 6 la_data_in[41]
port 36 nsew signal input
rlabel metal2 s 328642 0 328698 800 6 la_data_in[42]
port 37 nsew signal input
rlabel metal2 s 332874 0 332930 800 6 la_data_in[43]
port 38 nsew signal input
rlabel metal2 s 337106 0 337162 800 6 la_data_in[44]
port 39 nsew signal input
rlabel metal2 s 341338 0 341394 800 6 la_data_in[45]
port 40 nsew signal input
rlabel metal2 s 345570 0 345626 800 6 la_data_in[46]
port 41 nsew signal input
rlabel metal2 s 349802 0 349858 800 6 la_data_in[47]
port 42 nsew signal input
rlabel metal2 s 354034 0 354090 800 6 la_data_in[48]
port 43 nsew signal input
rlabel metal2 s 358266 0 358322 800 6 la_data_in[49]
port 44 nsew signal input
rlabel metal2 s 45098 0 45154 800 6 la_data_in[4]
port 45 nsew signal input
rlabel metal2 s 362498 0 362554 800 6 la_data_in[50]
port 46 nsew signal input
rlabel metal2 s 366730 0 366786 800 6 la_data_in[51]
port 47 nsew signal input
rlabel metal2 s 370962 0 371018 800 6 la_data_in[52]
port 48 nsew signal input
rlabel metal2 s 375194 0 375250 800 6 la_data_in[53]
port 49 nsew signal input
rlabel metal2 s 379426 0 379482 800 6 la_data_in[54]
port 50 nsew signal input
rlabel metal2 s 383658 0 383714 800 6 la_data_in[55]
port 51 nsew signal input
rlabel metal2 s 387890 0 387946 800 6 la_data_in[56]
port 52 nsew signal input
rlabel metal2 s 392122 0 392178 800 6 la_data_in[57]
port 53 nsew signal input
rlabel metal2 s 396354 0 396410 800 6 la_data_in[58]
port 54 nsew signal input
rlabel metal2 s 400586 0 400642 800 6 la_data_in[59]
port 55 nsew signal input
rlabel metal2 s 53562 0 53618 800 6 la_data_in[5]
port 56 nsew signal input
rlabel metal2 s 404818 0 404874 800 6 la_data_in[60]
port 57 nsew signal input
rlabel metal2 s 409050 0 409106 800 6 la_data_in[61]
port 58 nsew signal input
rlabel metal2 s 413282 0 413338 800 6 la_data_in[62]
port 59 nsew signal input
rlabel metal2 s 417514 0 417570 800 6 la_data_in[63]
port 60 nsew signal input
rlabel metal2 s 421746 0 421802 800 6 la_data_in[64]
port 61 nsew signal input
rlabel metal2 s 425978 0 426034 800 6 la_data_in[65]
port 62 nsew signal input
rlabel metal2 s 430210 0 430266 800 6 la_data_in[66]
port 63 nsew signal input
rlabel metal2 s 434442 0 434498 800 6 la_data_in[67]
port 64 nsew signal input
rlabel metal2 s 438674 0 438730 800 6 la_data_in[68]
port 65 nsew signal input
rlabel metal2 s 442906 0 442962 800 6 la_data_in[69]
port 66 nsew signal input
rlabel metal2 s 62026 0 62082 800 6 la_data_in[6]
port 67 nsew signal input
rlabel metal2 s 447138 0 447194 800 6 la_data_in[70]
port 68 nsew signal input
rlabel metal2 s 451370 0 451426 800 6 la_data_in[71]
port 69 nsew signal input
rlabel metal2 s 455602 0 455658 800 6 la_data_in[72]
port 70 nsew signal input
rlabel metal2 s 459834 0 459890 800 6 la_data_in[73]
port 71 nsew signal input
rlabel metal2 s 464066 0 464122 800 6 la_data_in[74]
port 72 nsew signal input
rlabel metal2 s 468298 0 468354 800 6 la_data_in[75]
port 73 nsew signal input
rlabel metal2 s 472530 0 472586 800 6 la_data_in[76]
port 74 nsew signal input
rlabel metal2 s 476762 0 476818 800 6 la_data_in[77]
port 75 nsew signal input
rlabel metal2 s 480994 0 481050 800 6 la_data_in[78]
port 76 nsew signal input
rlabel metal2 s 485226 0 485282 800 6 la_data_in[79]
port 77 nsew signal input
rlabel metal2 s 70490 0 70546 800 6 la_data_in[7]
port 78 nsew signal input
rlabel metal2 s 489458 0 489514 800 6 la_data_in[80]
port 79 nsew signal input
rlabel metal2 s 493690 0 493746 800 6 la_data_in[81]
port 80 nsew signal input
rlabel metal2 s 497922 0 497978 800 6 la_data_in[82]
port 81 nsew signal input
rlabel metal2 s 502154 0 502210 800 6 la_data_in[83]
port 82 nsew signal input
rlabel metal2 s 506386 0 506442 800 6 la_data_in[84]
port 83 nsew signal input
rlabel metal2 s 510618 0 510674 800 6 la_data_in[85]
port 84 nsew signal input
rlabel metal2 s 514850 0 514906 800 6 la_data_in[86]
port 85 nsew signal input
rlabel metal2 s 519082 0 519138 800 6 la_data_in[87]
port 86 nsew signal input
rlabel metal2 s 523314 0 523370 800 6 la_data_in[88]
port 87 nsew signal input
rlabel metal2 s 527546 0 527602 800 6 la_data_in[89]
port 88 nsew signal input
rlabel metal2 s 78954 0 79010 800 6 la_data_in[8]
port 89 nsew signal input
rlabel metal2 s 531778 0 531834 800 6 la_data_in[90]
port 90 nsew signal input
rlabel metal2 s 536010 0 536066 800 6 la_data_in[91]
port 91 nsew signal input
rlabel metal2 s 540242 0 540298 800 6 la_data_in[92]
port 92 nsew signal input
rlabel metal2 s 544474 0 544530 800 6 la_data_in[93]
port 93 nsew signal input
rlabel metal2 s 548706 0 548762 800 6 la_data_in[94]
port 94 nsew signal input
rlabel metal2 s 552938 0 552994 800 6 la_data_in[95]
port 95 nsew signal input
rlabel metal2 s 87418 0 87474 800 6 la_data_in[9]
port 96 nsew signal input
rlabel metal2 s 15474 0 15530 800 6 la_data_out[0]
port 97 nsew signal output
rlabel metal2 s 100114 0 100170 800 6 la_data_out[10]
port 98 nsew signal output
rlabel metal2 s 108578 0 108634 800 6 la_data_out[11]
port 99 nsew signal output
rlabel metal2 s 117042 0 117098 800 6 la_data_out[12]
port 100 nsew signal output
rlabel metal2 s 125506 0 125562 800 6 la_data_out[13]
port 101 nsew signal output
rlabel metal2 s 133970 0 134026 800 6 la_data_out[14]
port 102 nsew signal output
rlabel metal2 s 142434 0 142490 800 6 la_data_out[15]
port 103 nsew signal output
rlabel metal2 s 150898 0 150954 800 6 la_data_out[16]
port 104 nsew signal output
rlabel metal2 s 159362 0 159418 800 6 la_data_out[17]
port 105 nsew signal output
rlabel metal2 s 167826 0 167882 800 6 la_data_out[18]
port 106 nsew signal output
rlabel metal2 s 176290 0 176346 800 6 la_data_out[19]
port 107 nsew signal output
rlabel metal2 s 23938 0 23994 800 6 la_data_out[1]
port 108 nsew signal output
rlabel metal2 s 184754 0 184810 800 6 la_data_out[20]
port 109 nsew signal output
rlabel metal2 s 193218 0 193274 800 6 la_data_out[21]
port 110 nsew signal output
rlabel metal2 s 201682 0 201738 800 6 la_data_out[22]
port 111 nsew signal output
rlabel metal2 s 210146 0 210202 800 6 la_data_out[23]
port 112 nsew signal output
rlabel metal2 s 218610 0 218666 800 6 la_data_out[24]
port 113 nsew signal output
rlabel metal2 s 227074 0 227130 800 6 la_data_out[25]
port 114 nsew signal output
rlabel metal2 s 235538 0 235594 800 6 la_data_out[26]
port 115 nsew signal output
rlabel metal2 s 244002 0 244058 800 6 la_data_out[27]
port 116 nsew signal output
rlabel metal2 s 252466 0 252522 800 6 la_data_out[28]
port 117 nsew signal output
rlabel metal2 s 260930 0 260986 800 6 la_data_out[29]
port 118 nsew signal output
rlabel metal2 s 32402 0 32458 800 6 la_data_out[2]
port 119 nsew signal output
rlabel metal2 s 269394 0 269450 800 6 la_data_out[30]
port 120 nsew signal output
rlabel metal2 s 277858 0 277914 800 6 la_data_out[31]
port 121 nsew signal output
rlabel metal2 s 286322 0 286378 800 6 la_data_out[32]
port 122 nsew signal output
rlabel metal2 s 40866 0 40922 800 6 la_data_out[3]
port 123 nsew signal output
rlabel metal2 s 49330 0 49386 800 6 la_data_out[4]
port 124 nsew signal output
rlabel metal2 s 57794 0 57850 800 6 la_data_out[5]
port 125 nsew signal output
rlabel metal2 s 66258 0 66314 800 6 la_data_out[6]
port 126 nsew signal output
rlabel metal2 s 74722 0 74778 800 6 la_data_out[7]
port 127 nsew signal output
rlabel metal2 s 83186 0 83242 800 6 la_data_out[8]
port 128 nsew signal output
rlabel metal2 s 91650 0 91706 800 6 la_data_out[9]
port 129 nsew signal output
rlabel metal4 s 4208 2128 4528 349840 6 vccd1
port 130 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 349840 6 vccd1
port 130 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 349840 6 vccd1
port 130 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 349840 6 vccd1
port 130 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 349840 6 vccd1
port 130 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 349840 6 vccd1
port 130 nsew power bidirectional
rlabel metal4 s 188528 2128 188848 349840 6 vccd1
port 130 nsew power bidirectional
rlabel metal4 s 219248 2128 219568 349840 6 vccd1
port 130 nsew power bidirectional
rlabel metal4 s 249968 2128 250288 349840 6 vccd1
port 130 nsew power bidirectional
rlabel metal4 s 280688 2128 281008 349840 6 vccd1
port 130 nsew power bidirectional
rlabel metal4 s 311408 2128 311728 349840 6 vccd1
port 130 nsew power bidirectional
rlabel metal4 s 342128 2128 342448 349840 6 vccd1
port 130 nsew power bidirectional
rlabel metal4 s 372848 2128 373168 349840 6 vccd1
port 130 nsew power bidirectional
rlabel metal4 s 403568 2128 403888 349840 6 vccd1
port 130 nsew power bidirectional
rlabel metal4 s 434288 2128 434608 349840 6 vccd1
port 130 nsew power bidirectional
rlabel metal4 s 465008 2128 465328 349840 6 vccd1
port 130 nsew power bidirectional
rlabel metal4 s 495728 2128 496048 349840 6 vccd1
port 130 nsew power bidirectional
rlabel metal4 s 526448 2128 526768 349840 6 vccd1
port 130 nsew power bidirectional
rlabel metal4 s 557168 2128 557488 349840 6 vccd1
port 130 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 349840 6 vssd1
port 131 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 349840 6 vssd1
port 131 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 349840 6 vssd1
port 131 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 349840 6 vssd1
port 131 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 349840 6 vssd1
port 131 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 349840 6 vssd1
port 131 nsew ground bidirectional
rlabel metal4 s 203888 2128 204208 349840 6 vssd1
port 131 nsew ground bidirectional
rlabel metal4 s 234608 2128 234928 349840 6 vssd1
port 131 nsew ground bidirectional
rlabel metal4 s 265328 2128 265648 349840 6 vssd1
port 131 nsew ground bidirectional
rlabel metal4 s 296048 2128 296368 349840 6 vssd1
port 131 nsew ground bidirectional
rlabel metal4 s 326768 2128 327088 349840 6 vssd1
port 131 nsew ground bidirectional
rlabel metal4 s 357488 2128 357808 349840 6 vssd1
port 131 nsew ground bidirectional
rlabel metal4 s 388208 2128 388528 349840 6 vssd1
port 131 nsew ground bidirectional
rlabel metal4 s 418928 2128 419248 349840 6 vssd1
port 131 nsew ground bidirectional
rlabel metal4 s 449648 2128 449968 349840 6 vssd1
port 131 nsew ground bidirectional
rlabel metal4 s 480368 2128 480688 349840 6 vssd1
port 131 nsew ground bidirectional
rlabel metal4 s 511088 2128 511408 349840 6 vssd1
port 131 nsew ground bidirectional
rlabel metal4 s 541808 2128 542128 349840 6 vssd1
port 131 nsew ground bidirectional
rlabel metal2 s 7010 0 7066 800 6 wb_clk_i
port 132 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 560000 352000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 63396456
string GDS_FILE /home/mark/efabless_2023/caravel_template/openlane/user_proj_example/runs/23_09_01_13_33/results/signoff/user_proj_example.magic.gds
string GDS_START 978812
<< end >>

