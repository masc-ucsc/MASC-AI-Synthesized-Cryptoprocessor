module __masc__execute(
  input wire clk,
  input wire [31:0] instruction,
  input wire [31:0] rs1,
  input wire [31:0] rs2,
  output wire [32:0] out
);
  // ===== Pipe stage 0:

  // Registers for pipe stage 0:
  reg [31:0] p0_instruction;
  reg [31:0] p0_rs1;
  reg [31:0] p0_rs2;
  always_ff @ (posedge clk) begin
    p0_instruction <= instruction;
    p0_rs1 <= rs1;
    p0_rs2 <= rs2;
  end

  // ===== Pipe stage 1:
  wire p1_literal_11276_comb;
  wire [4:0] p1_bit_slice_11277_comb;
  wire [5:0] p1_literal_11278_comb;
  wire [5:0] p1_concat_11279_comb;
  wire [31:0] p1_literal_11280_comb;
  wire p1_rotation_1__8_comb;
  wire [30:0] p1_rotation_1__7_comb;
  wire [7:0] p1_byte0__1_comb;
  wire [23:0] p1_rotation_2__7_comb;
  wire [27:0] p1_rotation_1__12_comb;
  wire [3:0] p1_rotation_1__11_comb;
  wire [1:0] p1_rotation_2__12_comb;
  wire [29:0] p1_rotation_2__11_comb;
  wire [31:0] p1_literal_11289_comb;
  wire [31:0] p1_literal_11290_comb;
  wire [31:0] p1_literal_11291_comb;
  wire [31:0] p1_literal_11292_comb;
  wire [5:0] p1_sub_11293_comb;
  wire [31:0] p1_sub_11294_comb;
  wire [6:0] p1_literal_11295_comb;
  wire [24:0] p1_rotation_3__4_comb;
  wire [31:0] p1_rotation_1__1_comb;
  wire [31:0] p1_rotation_2__1_comb;
  wire [31:0] p1_rotation_1__2_comb;
  wire [31:0] p1_rotation_2__2_comb;
  wire [6:0] p1_rotation_3__5_comb;
  wire [1:0] p1_bit_slice_11302_comb;
  wire [1:0] p1_bit_slice_11303_comb;
  wire [20:0] p1_bit_slice_11304_comb;
  wire [20:0] p1_bit_slice_11305_comb;
  wire [20:0] p1_bit_slice_11306_comb;
  wire [1:0] p1_bit_slice_11307_comb;
  wire [1:0] p1_bit_slice_11308_comb;
  wire [10:0] p1_bit_slice_11309_comb;
  wire [10:0] p1_bit_slice_11310_comb;
  wire [10:0] p1_bit_slice_11311_comb;
  wire [2:0] p1_bit_slice_11312_comb;
  wire [2:0] p1_bit_slice_11313_comb;
  wire [10:0] p1_bit_slice_11314_comb;
  wire [5:0] p1_rotation_1__14_comb;
  wire [5:0] p1_bit_slice_11316_comb;
  wire [5:0] p1_bit_slice_11317_comb;
  wire [4:0] p1_bit_slice_11318_comb;
  wire [4:0] p1_bit_slice_11319_comb;
  wire [4:0] p1_bit_slice_11320_comb;
  wire [5:0] p1_bit_slice_11321_comb;
  wire [5:0] p1_rotation_2__18_comb;
  wire [9:0] p1_bit_slice_11323_comb;
  wire [9:0] p1_bit_slice_11324_comb;
  wire [5:0] p1_bit_slice_11325_comb;
  wire [5:0] p1_bit_slice_11326_comb;
  wire [12:0] p1_bit_slice_11327_comb;
  wire [12:0] p1_bit_slice_11328_comb;
  wire [12:0] p1_rotation_1__19_comb;
  wire [31:0] p1_literal_11330_comb;
  wire [8:0] p1_bit_slice_11331_comb;
  wire [8:0] p1_bit_slice_11332_comb;
  wire [8:0] p1_bit_slice_11333_comb;
  wire [13:0] p1_bit_slice_11334_comb;
  wire [13:0] p1_rotate_18__1_comb;
  wire [13:0] p1_bit_slice_11336_comb;
  wire [3:0] p1_bit_slice_11337_comb;
  wire [3:0] p1_bit_slice_11338_comb;
  wire [9:0] p1_bit_slice_11339_comb;
  wire [9:0] p1_bit_slice_11340_comb;
  wire [6:0] p1_bit_slice_11341_comb;
  wire [6:0] p1_rotation_3__6_comb;
  wire [6:0] p1_bit_slice_11343_comb;
  wire [9:0] p1_bit_slice_11344_comb;
  wire [9:0] p1_bit_slice_11345_comb;
  wire [9:0] p1_rot_c__1_comb;
  wire [13:0] p1_bit_slice_11347_comb;
  wire [13:0] p1_bit_slice_11348_comb;
  wire [13:0] p1_bit_slice_11349_comb;
  wire [13:0] p1_bit_slice_11350_comb;
  wire [12:0] p1_bit_slice_11351_comb;
  wire [3:0] p1_bit_slice_11352_comb;
  wire [3:0] p1_bit_slice_11353_comb;
  wire [6:0] p1_bit_slice_11354_comb;
  wire [6:0] p1_bit_slice_11355_comb;
  wire [2:0] p1_bit_slice_11356_comb;
  wire [2:0] p1_rotation_2__19_comb;
  wire [2:0] p1_bit_slice_11358_comb;
  wire p1_eq_11359_comb;
  wire p1_eq_11360_comb;
  wire [31:0] p1_literal_11361_comb;
  wire [31:0] p1_literal_11362_comb;
  wire [31:0] p1_literal_11363_comb;
  wire [31:0] p1_literal_11364_comb;
  wire [31:0] p1_literal_11365_comb;
  wire [31:0] p1_literal_11366_comb;
  wire [31:0] p1_literal_11367_comb;
  wire [31:0] p1_literal_11368_comb;
  wire [31:0] p1_literal_11369_comb;
  wire [31:0] p1_literal_11370_comb;
  wire p1_eq_11371_comb;
  wire p1_eq_11372_comb;
  wire [31:0] p1_literal_11373_comb;
  wire [31:0] p1_literal_11374_comb;
  wire [31:0] p1_literal_11375_comb;
  wire [31:0] p1_literal_11376_comb;
  wire [31:0] p1_literal_11377_comb;
  wire [31:0] p1_literal_11378_comb;
  wire [31:0] p1_literal_11379_comb;
  wire [31:0] p1_shrl_11380_comb;
  wire [31:0] p1_shll_11381_comb;
  wire [31:0] p1_shll_11382_comb;
  wire [31:0] p1_shrl_11383_comb;
  wire [31:0] p1_shrl_11384_comb;
  wire [31:0] p1_shll_11385_comb;
  wire [31:0] p1_not_11386_comb;
  wire [31:0] p1_xor_11387_comb;
  wire [31:0] p1_shift_1_comb;
  wire [31:0] p1_combined_1_comb;
  wire [31:0] p1_combined_2_comb;
  wire [8:0] p1_bit_slice_11391_comb;
  wire [8:0] p1_bit_slice_11392_comb;
  wire [8:0] p1_rotation_3__9_comb;
  wire [31:0] p1_combined_1__1_comb;
  wire [31:0] p1_combined_2__1_comb;
  wire [31:0] p1_rotation_3__1_comb;
  wire [1:0] p1_result__39_comb;
  wire [4:0] p1_bit_slice_11398_comb;
  wire [20:0] p1_result__37_comb;
  wire [1:0] p1_xor_11400_comb;
  wire [10:0] p1_xor_11401_comb;
  wire [2:0] p1_xor_11402_comb;
  wire [3:0] p1_bit_slice_11403_comb;
  wire [10:0] p1_xor_11404_comb;
  wire [5:0] p1_xor_11405_comb;
  wire [4:0] p1_xor_11406_comb;
  wire [5:0] p1_result__47_comb;
  wire [9:0] p1_result__46_comb;
  wire [5:0] p1_xor_11409_comb;
  wire [12:0] p1_xor_11410_comb;
  wire p1_eq_11411_comb;
  wire [8:0] p1_xor_11412_comb;
  wire [13:0] p1_xor_11413_comb;
  wire [4:0] p1_bit_slice_11414_comb;
  wire [4:0] p1_bit_slice_11415_comb;
  wire [3:0] p1_result__41_comb;
  wire [9:0] p1_xor_11417_comb;
  wire [6:0] p1_xor_11418_comb;
  wire [6:0] p1_result__45_comb;
  wire [9:0] p1_xor_11420_comb;
  wire [13:0] p1_xor_11421_comb;
  wire [13:0] p1_result__40_comb;
  wire [9:0] p1_xor_11423_comb;
  wire [1:0] p1_bit_slice_11424_comb;
  wire [1:0] p1_bit_slice_11425_comb;
  wire [12:0] p1_xor_11426_comb;
  wire [8:0] p1_bit_slice_11427_comb;
  wire [8:0] p1_bit_slice_11428_comb;
  wire [3:0] p1_result__36_comb;
  wire [6:0] p1_xor_11430_comb;
  wire [2:0] p1_xor_11431_comb;
  wire p1_or_11432_comb;
  wire p1_eq_11433_comb;
  wire p1_eq_11434_comb;
  wire p1_eq_11435_comb;
  wire p1_eq_11436_comb;
  wire p1_eq_11437_comb;
  wire p1_eq_11438_comb;
  wire p1_eq_11439_comb;
  wire p1_eq_11440_comb;
  wire p1_eq_11441_comb;
  wire p1_eq_11442_comb;
  wire p1_or_11443_comb;
  wire p1_eq_11444_comb;
  wire p1_eq_11445_comb;
  wire p1_eq_11446_comb;
  wire p1_eq_11447_comb;
  wire p1_eq_11448_comb;
  wire p1_eq_11449_comb;
  wire p1_eq_11450_comb;
  wire [31:0] p1_or_11451_comb;
  wire [31:0] p1_or_11452_comb;
  wire [31:0] p1_or_11453_comb;
  wire [31:0] p1_nor_11454_comb;
  wire [31:0] p1_nand_11455_comb;
  wire [31:0] p1_not_11456_comb;
  wire [31:0] p1_xor_11457_comb;
  wire [8:0] p1_result__43_comb;
  wire [31:0] p1_xor_11459_comb;
  wire p1_result__23_comb;
  wire p1_result__25_comb;
  wire p1_result__27_comb;
  wire p1_result__29_comb;
  wire p1_result__31_comb;
  wire p1_result__33_comb;
  wire p1_result__35_comb;
  wire p1_result__34_comb;
  wire p1_result__32_comb;
  wire p1_result__30_comb;
  wire p1_result__28_comb;
  wire p1_result__19_comb;
  wire p1_result__15_comb;
  wire p1_result__11_comb;
  wire p1_result__7_comb;
  wire p1_bit_slice_11475_comb;
  wire [4:0] p1_result__38_comb;
  wire p1_bit_slice_11477_comb;
  wire p1_bit_slice_11478_comb;
  wire [5:0] p1_bit_slice_11479_comb;
  wire [1:0] p1_bit_slice_11480_comb;
  wire [3:0] p1_xor_11481_comb;
  wire p1_bit_slice_11482_comb;
  wire [4:0] p1_bit_slice_11483_comb;
  wire [1:0] p1_bit_slice_11484_comb;
  wire [4:0] p1_bit_slice_11485_comb;
  wire [1:0] p1_bit_slice_11486_comb;
  wire [4:0] p1_bit_slice_11487_comb;
  wire [1:0] p1_bit_slice_11488_comb;
  wire p1_or_11489_comb;
  wire p1_result__9_comb;
  wire p1_result__13_comb;
  wire p1_result__17_comb;
  wire p1_result__26_comb;
  wire p1_result__24_comb;
  wire p1_result__22_comb;
  wire p1_result__21_comb;
  wire p1_result__18_comb;
  wire p1_result__14_comb;
  wire p1_result__10_comb;
  wire [3:0] p1_bit_slice_11500_comb;
  wire [1:0] p1_bit_slice_11501_comb;
  wire [1:0] p1_bit_slice_11502_comb;
  wire [3:0] p1_bit_slice_11503_comb;
  wire [4:0] p1_result__42_comb;
  wire p1_bit_slice_11505_comb;
  wire p1_bit_slice_11506_comb;
  wire [4:0] p1_bit_slice_11507_comb;
  wire p1_or_11508_comb;
  wire p1_bit_slice_11509_comb;
  wire p1_literal_11510_comb;
  wire p1_bit_slice_11511_comb;
  wire p1_result__20_comb;
  wire p1_result__6_comb;
  wire p1_bit_slice_11514_comb;
  wire p1_bit_slice_11515_comb;
  wire p1_result__16_comb;
  wire [4:0] p1_bit_slice_11517_comb;
  wire p1_bit_slice_11518_comb;
  wire p1_bit_slice_11519_comb;
  wire [4:0] p1_bit_slice_11520_comb;
  wire p1_bit_slice_11521_comb;
  wire [4:0] p1_bit_slice_11522_comb;
  wire [1:0] p1_bit_slice_11523_comb;
  wire [3:0] p1_bit_slice_11524_comb;
  wire [1:0] p1_xor_11525_comb;
  wire [3:0] p1_bit_slice_11526_comb;
  wire [8:0] p1_result__44_comb;
  wire p1_result__8_comb;
  wire p1_result__12_comb;
  wire p1_result__5_comb;
  wire [3:0] p1_bit_slice_11531_comb;
  wire [2:0] p1_bit_slice_11532_comb;
  wire p1_bit_slice_11533_comb;
  wire [5:0] p1_bit_slice_11534_comb;
  wire [4:0] p1_bit_slice_11535_comb;
  wire [1:0] p1_bit_slice_11536_comb;
  wire p1_or_11537_comb;
  wire [19:0] p1_concat_11538_comb;
  wire p1_bit_slice_11539_comb;
  wire p1_bit_slice_11540_comb;
  wire p1_bit_slice_11541_comb;
  wire p1_bit_slice_11542_comb;
  wire p1_bit_slice_11543_comb;
  wire p1_bit_slice_11544_comb;
  wire p1_bit_slice_11545_comb;
  wire p1_bit_slice_11546_comb;
  wire p1_bit_slice_11547_comb;
  wire p1_bit_slice_11548_comb;
  wire p1_bit_slice_11549_comb;
  wire p1_bit_slice_11550_comb;
  wire p1_bit_slice_11551_comb;
  wire p1_bit_slice_11552_comb;
  wire p1_bit_slice_11553_comb;
  wire p1_bit_slice_11554_comb;
  wire p1_bit_slice_11555_comb;
  wire [20:0] p1_concat_11556_comb;
  wire [6:0] p1_bit_slice_11557_comb;
  wire [6:0] p1_bit_slice_11558_comb;
  wire [6:0] p1_bit_slice_11559_comb;
  wire [6:0] p1_bit_slice_11560_comb;
  wire [6:0] p1_bit_slice_11561_comb;
  wire [6:0] p1_bit_slice_11562_comb;
  wire [6:0] p1_bit_slice_11563_comb;
  wire [6:0] p1_concat_11564_comb;
  wire [6:0] p1_concat_11565_comb;
  wire [6:0] p1_concat_11566_comb;
  wire [6:0] p1_concat_11567_comb;
  wire [6:0] p1_concat_11568_comb;
  wire [6:0] p1_bit_slice_11569_comb;
  wire [6:0] p1_concat_11570_comb;
  wire [6:0] p1_concat_11571_comb;
  wire [6:0] p1_bit_slice_11572_comb;
  wire [6:0] p1_bit_slice_11573_comb;
  wire [6:0] p1_concat_11574_comb;
  wire [6:0] p1_concat_11575_comb;
  wire [6:0] p1_bit_slice_11576_comb;
  wire [19:0] p1_concat_11577_comb;
  wire p1_bit_slice_11578_comb;
  wire p1_bit_slice_11579_comb;
  wire p1_bit_slice_11580_comb;
  wire p1_bit_slice_11581_comb;
  wire p1_bit_slice_11582_comb;
  wire p1_bit_slice_11583_comb;
  wire p1_bit_slice_11584_comb;
  wire p1_bit_slice_11585_comb;
  wire p1_bit_slice_11586_comb;
  wire p1_bit_slice_11587_comb;
  wire p1_bit_slice_11588_comb;
  wire p1_bit_slice_11589_comb;
  wire p1_bit_slice_11590_comb;
  wire p1_bit_slice_11591_comb;
  wire p1_bit_slice_11592_comb;
  wire p1_bit_slice_11593_comb;
  wire [5:0] p1_bit_slice_11594_comb;
  wire [5:0] p1_bit_slice_11595_comb;
  wire [5:0] p1_bit_slice_11596_comb;
  wire [5:0] p1_bit_slice_11597_comb;
  wire [5:0] p1_bit_slice_11598_comb;
  wire [5:0] p1_bit_slice_11599_comb;
  wire [5:0] p1_bit_slice_11600_comb;
  wire [5:0] p1_concat_11601_comb;
  wire [5:0] p1_bit_slice_11602_comb;
  wire [5:0] p1_concat_11603_comb;
  wire [5:0] p1_concat_11604_comb;
  wire [5:0] p1_bit_slice_11605_comb;
  wire [5:0] p1_concat_11606_comb;
  wire [5:0] p1_bit_slice_11607_comb;
  wire [5:0] p1_bit_slice_11608_comb;
  wire [5:0] p1_concat_11609_comb;
  wire [5:0] p1_concat_11610_comb;
  wire [5:0] p1_bit_slice_11611_comb;
  wire [5:0] p1_bit_slice_11612_comb;
  wire [5:0] p1_bit_slice_11613_comb;
  wire [5:0] p1_concat_11614_comb;
  wire [20:0] p1_concat_11615_comb;
  wire [1:0] p1_bit_slice_11616_comb;
  wire [1:0] p1_bit_slice_11617_comb;
  wire [1:0] p1_bit_slice_11618_comb;
  wire [1:0] p1_bit_slice_11619_comb;
  wire [1:0] p1_bit_slice_11620_comb;
  wire [1:0] p1_bit_slice_11621_comb;
  wire [1:0] p1_concat_11622_comb;
  wire [1:0] p1_concat_11623_comb;
  wire [1:0] p1_concat_11624_comb;
  wire [1:0] p1_concat_11625_comb;
  wire [1:0] p1_concat_11626_comb;
  wire [1:0] p1_bit_slice_11627_comb;
  wire [1:0] p1_bit_slice_11628_comb;
  wire [1:0] p1_bit_slice_11629_comb;
  wire [1:0] p1_bit_slice_11630_comb;
  wire [1:0] p1_bit_slice_11631_comb;
  wire [1:0] p1_bit_slice_11632_comb;
  wire [1:0] p1_bit_slice_11633_comb;
  wire [1:0] p1_concat_11634_comb;
  wire [1:0] p1_bit_slice_11635_comb;
  wire [1:0] p1_bit_slice_11636_comb;
  wire [21:0] p1_concat_11637_comb;
  wire [5:0] p1_bit_slice_11638_comb;
  wire [5:0] p1_bit_slice_11639_comb;
  wire [5:0] p1_bit_slice_11640_comb;
  wire [5:0] p1_bit_slice_11641_comb;
  wire [5:0] p1_bit_slice_11642_comb;
  wire [5:0] p1_bit_slice_11643_comb;
  wire [5:0] p1_concat_11644_comb;
  wire [5:0] p1_bit_slice_11645_comb;
  wire [5:0] p1_concat_11646_comb;
  wire [5:0] p1_concat_11647_comb;
  wire [5:0] p1_bit_slice_11648_comb;
  wire [5:0] p1_concat_11649_comb;
  wire [5:0] p1_bit_slice_11650_comb;
  wire [5:0] p1_concat_11651_comb;
  wire [5:0] p1_bit_slice_11652_comb;
  wire [5:0] p1_concat_11653_comb;
  wire [5:0] p1_bit_slice_11654_comb;
  wire [5:0] p1_bit_slice_11655_comb;
  wire [5:0] p1_concat_11656_comb;
  wire [5:0] p1_concat_11657_comb;
  wire [20:0] p1_concat_11658_comb;
  wire p1_bit_slice_11659_comb;
  wire p1_bit_slice_11660_comb;
  wire p1_bit_slice_11661_comb;
  wire p1_bit_slice_11662_comb;
  wire p1_bit_slice_11663_comb;
  wire p1_bit_slice_11664_comb;
  wire p1_bit_slice_11665_comb;
  wire p1_bit_slice_11666_comb;
  wire p1_bit_slice_11667_comb;
  wire p1_bit_slice_11668_comb;
  wire p1_bit_slice_11669_comb;
  wire p1_bit_slice_11670_comb;
  wire p1_bit_slice_11671_comb;
  wire p1_bit_slice_11672_comb;
  wire p1_bit_slice_11673_comb;
  wire p1_bit_slice_11674_comb;
  wire [20:0] p1_concat_11675_comb;
  wire [6:0] p1_bit_slice_11676_comb;
  wire [6:0] p1_bit_slice_11677_comb;
  wire [6:0] p1_bit_slice_11678_comb;
  wire [6:0] p1_bit_slice_11679_comb;
  wire [6:0] p1_bit_slice_11680_comb;
  wire [6:0] p1_bit_slice_11681_comb;
  wire [6:0] p1_bit_slice_11682_comb;
  wire [6:0] p1_concat_11683_comb;
  wire [6:0] p1_concat_11684_comb;
  wire [6:0] p1_concat_11685_comb;
  wire [6:0] p1_concat_11686_comb;
  wire [6:0] p1_bit_slice_11687_comb;
  wire [6:0] p1_bit_slice_11688_comb;
  wire [6:0] p1_bit_slice_11689_comb;
  wire [6:0] p1_concat_11690_comb;
  wire [6:0] p1_bit_slice_11691_comb;
  wire [6:0] p1_bit_slice_11692_comb;
  wire [6:0] p1_bit_slice_11693_comb;
  wire [6:0] p1_concat_11694_comb;
  wire [6:0] p1_bit_slice_11695_comb;
  wire [18:0] p1_concat_11696_comb;
  wire p1_bit_slice_11697_comb;
  wire p1_bit_slice_11698_comb;
  wire p1_bit_slice_11699_comb;
  wire p1_bit_slice_11700_comb;
  wire p1_bit_slice_11701_comb;
  wire p1_bit_slice_11702_comb;
  wire p1_bit_slice_11703_comb;
  wire p1_bit_slice_11704_comb;
  wire p1_bit_slice_11705_comb;
  wire p1_bit_slice_11706_comb;
  wire p1_bit_slice_11707_comb;
  wire p1_bit_slice_11708_comb;
  wire p1_bit_slice_11709_comb;
  wire p1_bit_slice_11710_comb;
  wire p1_bit_slice_11711_comb;
  wire p1_bit_slice_11712_comb;
  wire p1_one_hot_sel_11713_comb;
  wire [6:0] p1_one_hot_sel_11714_comb;
  wire p1_one_hot_sel_11715_comb;
  wire [5:0] p1_one_hot_sel_11716_comb;
  wire [1:0] p1_one_hot_sel_11717_comb;
  wire [5:0] p1_one_hot_sel_11718_comb;
  wire p1_one_hot_sel_11719_comb;
  wire [6:0] p1_one_hot_sel_11720_comb;
  wire p1_one_hot_sel_11721_comb;
  wire [31:0] p1_literal_11722_comb;
  wire [31:0] p1_concat_11723_comb;
  wire p1_ult_11724_comb;
  wire [32:0] p1_tuple_11725_comb;
  assign p1_literal_11276_comb = 1'h0;
  assign p1_bit_slice_11277_comb = p0_rs2[4:0];
  assign p1_literal_11278_comb = 6'h20;
  assign p1_concat_11279_comb = {p1_literal_11276_comb, p1_bit_slice_11277_comb};
  assign p1_literal_11280_comb = 32'h0000_0020;
  assign p1_rotation_1__8_comb = p0_rs1[0];
  assign p1_rotation_1__7_comb = p0_rs1[31:1];
  assign p1_byte0__1_comb = p0_rs1[7:0];
  assign p1_rotation_2__7_comb = p0_rs1[31:8];
  assign p1_rotation_1__12_comb = p0_rs1[27:0];
  assign p1_rotation_1__11_comb = p0_rs1[31:28];
  assign p1_rotation_2__12_comb = p0_rs1[1:0];
  assign p1_rotation_2__11_comb = p0_rs1[31:2];
  assign p1_literal_11289_comb = 32'h0000_0006;
  assign p1_literal_11290_comb = 32'h0000_0007;
  assign p1_literal_11291_comb = 32'h0000_000a;
  assign p1_literal_11292_comb = 32'h0000_000b;
  assign p1_sub_11293_comb = p1_literal_11278_comb - p1_concat_11279_comb;
  assign p1_sub_11294_comb = p1_literal_11280_comb - p0_rs2;
  assign p1_literal_11295_comb = 7'h00;
  assign p1_rotation_3__4_comb = p0_rs1[31:7];
  assign p1_rotation_1__1_comb = {p1_rotation_1__8_comb, p1_rotation_1__7_comb};
  assign p1_rotation_2__1_comb = {p1_byte0__1_comb, p1_rotation_2__7_comb};
  assign p1_rotation_1__2_comb = {p1_rotation_1__12_comb, p1_rotation_1__11_comb};
  assign p1_rotation_2__2_comb = {p1_rotation_2__12_comb, p1_rotation_2__11_comb};
  assign p1_rotation_3__5_comb = p0_rs1[6:0];
  assign p1_bit_slice_11302_comb = p0_rs1[27:26];
  assign p1_bit_slice_11303_comb = p0_rs1[6:5];
  assign p1_bit_slice_11304_comb = p0_rs1[20:0];
  assign p1_bit_slice_11305_comb = p0_rs1[26:6];
  assign p1_bit_slice_11306_comb = p0_rs1[31:11];
  assign p1_bit_slice_11307_comb = p0_rs1[12:11];
  assign p1_bit_slice_11308_comb = p0_rs1[21:20];
  assign p1_bit_slice_11309_comb = p0_rs1[31:21];
  assign p1_bit_slice_11310_comb = p0_rs1[10:0];
  assign p1_bit_slice_11311_comb = p0_rs1[19:9];
  assign p1_bit_slice_11312_comb = p0_rs1[6:4];
  assign p1_bit_slice_11313_comb = p0_rs1[17:15];
  assign p1_bit_slice_11314_comb = p0_rs1[27:17];
  assign p1_rotation_1__14_comb = p0_rs1[5:0];
  assign p1_bit_slice_11316_comb = p0_rs1[10:5];
  assign p1_bit_slice_11317_comb = p0_rs1[24:19];
  assign p1_bit_slice_11318_comb = p0_rs1[31:27];
  assign p1_bit_slice_11319_comb = p0_rs1[4:0];
  assign p1_bit_slice_11320_comb = p0_rs1[18:14];
  assign p1_bit_slice_11321_comb = p0_rs1[15:10];
  assign p1_rotation_2__18_comb = p0_rs2[5:0];
  assign p1_bit_slice_11323_comb = p0_rs1[9:0];
  assign p1_bit_slice_11324_comb = p0_rs2[31:22];
  assign p1_bit_slice_11325_comb = p0_rs1[18:13];
  assign p1_bit_slice_11326_comb = p0_rs1[28:23];
  assign p1_bit_slice_11327_comb = p0_rs1[12:0];
  assign p1_bit_slice_11328_comb = p0_rs1[22:10];
  assign p1_rotation_1__19_comb = p0_rs1[31:19];
  assign p1_literal_11330_comb = 32'h0000_0009;
  assign p1_bit_slice_11331_comb = p0_rs1[20:12];
  assign p1_bit_slice_11332_comb = p0_rs1[31:23];
  assign p1_bit_slice_11333_comb = p0_rs1[8:0];
  assign p1_bit_slice_11334_comb = p0_rs1[26:13];
  assign p1_rotate_18__1_comb = p0_rs1[31:18];
  assign p1_bit_slice_11336_comb = p0_rs1[13:0];
  assign p1_bit_slice_11337_comb = p0_rs1[3:0];
  assign p1_bit_slice_11338_comb = p0_rs2[26:23];
  assign p1_bit_slice_11339_comb = p0_rs1[16:7];
  assign p1_bit_slice_11340_comb = p0_rs1[18:9];
  assign p1_bit_slice_11341_comb = p0_rs1[8:2];
  assign p1_rotation_3__6_comb = p0_rs1[31:25];
  assign p1_bit_slice_11343_comb = p0_rs2[21:15];
  assign p1_bit_slice_11344_comb = p0_rs1[11:2];
  assign p1_bit_slice_11345_comb = p0_rs1[22:13];
  assign p1_rot_c__1_comb = p0_rs1[31:22];
  assign p1_bit_slice_11347_comb = p0_rs1[20:7];
  assign p1_bit_slice_11348_comb = p0_rs1[16:3];
  assign p1_bit_slice_11349_comb = p0_rs1[27:14];
  assign p1_bit_slice_11350_comb = p0_rs2[22:9];
  assign p1_bit_slice_11351_comb = p0_rs1[29:17];
  assign p1_bit_slice_11352_comb = p0_rs1[5:2];
  assign p1_bit_slice_11353_comb = p0_rs1[10:7];
  assign p1_bit_slice_11354_comb = p0_rs1[12:6];
  assign p1_bit_slice_11355_comb = p0_rs1[17:11];
  assign p1_bit_slice_11356_comb = p0_rs1[21:19];
  assign p1_rotation_2__19_comb = p0_rs1[31:29];
  assign p1_bit_slice_11358_comb = p0_rs1[8:6];
  assign p1_eq_11359_comb = p0_instruction == p1_literal_11289_comb;
  assign p1_eq_11360_comb = p0_instruction == p1_literal_11290_comb;
  assign p1_literal_11361_comb = 32'h0000_0015;
  assign p1_literal_11362_comb = 32'h0000_0014;
  assign p1_literal_11363_comb = 32'h0000_0013;
  assign p1_literal_11364_comb = 32'h0000_0012;
  assign p1_literal_11365_comb = 32'h0000_0011;
  assign p1_literal_11366_comb = 32'h0000_0010;
  assign p1_literal_11367_comb = 32'h0000_000f;
  assign p1_literal_11368_comb = 32'h0000_000e;
  assign p1_literal_11369_comb = 32'h0000_000d;
  assign p1_literal_11370_comb = 32'h0000_000c;
  assign p1_eq_11371_comb = p0_instruction == p1_literal_11291_comb;
  assign p1_eq_11372_comb = p0_instruction == p1_literal_11292_comb;
  assign p1_literal_11373_comb = 32'h0000_0008;
  assign p1_literal_11374_comb = 32'h0000_0005;
  assign p1_literal_11375_comb = 32'h0000_0004;
  assign p1_literal_11376_comb = 32'h0000_0003;
  assign p1_literal_11377_comb = 32'h0000_0002;
  assign p1_literal_11378_comb = 32'h0000_0001;
  assign p1_literal_11379_comb = 32'h0000_0000;
  assign p1_shrl_11380_comb = p0_rs1 >> p1_bit_slice_11277_comb;
  assign p1_shll_11381_comb = p1_sub_11293_comb >= 6'h20 ? 32'h0000_0000 : p0_rs1 << p1_sub_11293_comb;
  assign p1_shll_11382_comb = p0_rs1 << p1_bit_slice_11277_comb;
  assign p1_shrl_11383_comb = p1_sub_11293_comb >= 6'h20 ? 32'h0000_0000 : p0_rs1 >> p1_sub_11293_comb;
  assign p1_shrl_11384_comb = p0_rs2 >= 32'h0000_0020 ? 32'h0000_0000 : p0_rs1 >> p0_rs2;
  assign p1_shll_11385_comb = p1_sub_11294_comb >= 32'h0000_0020 ? 32'h0000_0000 : p0_rs1 << p1_sub_11294_comb;
  assign p1_not_11386_comb = ~p0_rs1;
  assign p1_xor_11387_comb = p0_rs1 ^ p0_rs2;
  assign p1_shift_1_comb = {p1_literal_11295_comb, p1_rotation_3__4_comb};
  assign p1_combined_1_comb = p1_rotation_1__1_comb & p0_rs2;
  assign p1_combined_2_comb = p1_rotation_2__1_comb | p0_rs2;
  assign p1_bit_slice_11391_comb = p0_rs1[13:5];
  assign p1_bit_slice_11392_comb = p0_rs1[17:9];
  assign p1_rotation_3__9_comb = p0_rs2[8:0];
  assign p1_combined_1__1_comb = p1_rotation_1__2_comb & p0_rs2;
  assign p1_combined_2__1_comb = p1_rotation_2__2_comb | p0_rs2;
  assign p1_rotation_3__1_comb = {p1_rotation_3__5_comb, p1_rotation_3__4_comb};
  assign p1_result__39_comb = p1_bit_slice_11302_comb ^ p1_rotation_2__12_comb ^ p1_bit_slice_11303_comb;
  assign p1_bit_slice_11398_comb = p0_rs1[25:21];
  assign p1_result__37_comb = p1_bit_slice_11304_comb ^ p1_bit_slice_11305_comb ^ p1_bit_slice_11306_comb;
  assign p1_xor_11400_comb = p1_rotation_2__12_comb ^ p1_bit_slice_11307_comb ^ p1_bit_slice_11308_comb;
  assign p1_xor_11401_comb = p1_bit_slice_11309_comb ^ p1_bit_slice_11310_comb ^ p1_bit_slice_11311_comb;
  assign p1_xor_11402_comb = p1_bit_slice_11312_comb ^ p1_bit_slice_11313_comb;
  assign p1_bit_slice_11403_comb = p0_rs1[14:11];
  assign p1_xor_11404_comb = p1_bit_slice_11309_comb ^ p1_bit_slice_11310_comb ^ p1_bit_slice_11314_comb;
  assign p1_xor_11405_comb = p1_rotation_1__14_comb ^ p1_bit_slice_11316_comb ^ p1_bit_slice_11317_comb;
  assign p1_xor_11406_comb = p1_bit_slice_11318_comb ^ p1_bit_slice_11319_comb ^ p1_bit_slice_11320_comb;
  assign p1_result__47_comb = p1_bit_slice_11321_comb ^ p1_rotation_2__18_comb;
  assign p1_result__46_comb = p1_bit_slice_11323_comb ^ p1_bit_slice_11324_comb;
  assign p1_xor_11409_comb = p1_bit_slice_11325_comb ^ p1_bit_slice_11326_comb;
  assign p1_xor_11410_comb = p1_bit_slice_11327_comb ^ p1_bit_slice_11328_comb ^ p1_rotation_1__19_comb;
  assign p1_eq_11411_comb = p0_instruction == p1_literal_11330_comb;
  assign p1_xor_11412_comb = p1_bit_slice_11331_comb ^ p1_bit_slice_11332_comb ^ p1_bit_slice_11333_comb;
  assign p1_xor_11413_comb = p1_bit_slice_11334_comb ^ p1_rotate_18__1_comb ^ p1_bit_slice_11336_comb;
  assign p1_bit_slice_11414_comb = p0_rs1[8:4];
  assign p1_bit_slice_11415_comb = p0_rs2[31:27];
  assign p1_result__41_comb = p1_rotation_1__11_comb ^ p1_bit_slice_11337_comb ^ p1_bit_slice_11338_comb;
  assign p1_xor_11417_comb = p1_bit_slice_11339_comb ^ p1_bit_slice_11340_comb;
  assign p1_xor_11418_comb = p1_rotation_3__5_comb ^ p1_bit_slice_11341_comb ^ p1_rotation_3__6_comb;
  assign p1_result__45_comb = p1_rotation_3__6_comb ^ p1_bit_slice_11343_comb;
  assign p1_xor_11420_comb = p1_bit_slice_11344_comb ^ p1_bit_slice_11345_comb ^ p1_rot_c__1_comb;
  assign p1_xor_11421_comb = p1_bit_slice_11347_comb ^ p1_rotate_18__1_comb ^ p1_bit_slice_11348_comb;
  assign p1_result__40_comb = p1_bit_slice_11349_comb ^ p1_rotate_18__1_comb ^ p1_bit_slice_11350_comb;
  assign p1_xor_11423_comb = p1_rot_c__1_comb ^ p1_bit_slice_11323_comb ^ p1_bit_slice_11340_comb;
  assign p1_bit_slice_11424_comb = p0_rs1[31:30];
  assign p1_bit_slice_11425_comb = p0_rs1[24:23];
  assign p1_xor_11426_comb = p1_bit_slice_11351_comb ^ p1_rotation_1__19_comb ^ p1_bit_slice_11328_comb;
  assign p1_bit_slice_11427_comb = p0_rs1[24:16];
  assign p1_bit_slice_11428_comb = p0_rs2[14:6];
  assign p1_result__36_comb = p1_rotation_1__11_comb ^ p1_bit_slice_11352_comb ^ p1_bit_slice_11353_comb;
  assign p1_xor_11430_comb = p1_bit_slice_11354_comb ^ p1_bit_slice_11355_comb ^ p1_rotation_3__6_comb;
  assign p1_xor_11431_comb = p1_bit_slice_11356_comb ^ p1_rotation_2__19_comb ^ p1_bit_slice_11358_comb;
  assign p1_or_11432_comb = p1_eq_11359_comb | p1_eq_11360_comb;
  assign p1_eq_11433_comb = p0_instruction == p1_literal_11361_comb;
  assign p1_eq_11434_comb = p0_instruction == p1_literal_11362_comb;
  assign p1_eq_11435_comb = p0_instruction == p1_literal_11363_comb;
  assign p1_eq_11436_comb = p0_instruction == p1_literal_11364_comb;
  assign p1_eq_11437_comb = p0_instruction == p1_literal_11365_comb;
  assign p1_eq_11438_comb = p0_instruction == p1_literal_11366_comb;
  assign p1_eq_11439_comb = p0_instruction == p1_literal_11367_comb;
  assign p1_eq_11440_comb = p0_instruction == p1_literal_11368_comb;
  assign p1_eq_11441_comb = p0_instruction == p1_literal_11369_comb;
  assign p1_eq_11442_comb = p0_instruction == p1_literal_11370_comb;
  assign p1_or_11443_comb = p1_eq_11371_comb | p1_eq_11372_comb;
  assign p1_eq_11444_comb = p0_instruction == p1_literal_11373_comb;
  assign p1_eq_11445_comb = p0_instruction == p1_literal_11374_comb;
  assign p1_eq_11446_comb = p0_instruction == p1_literal_11375_comb;
  assign p1_eq_11447_comb = p0_instruction == p1_literal_11376_comb;
  assign p1_eq_11448_comb = p0_instruction == p1_literal_11377_comb;
  assign p1_eq_11449_comb = p0_instruction == p1_literal_11378_comb;
  assign p1_eq_11450_comb = p0_instruction == p1_literal_11379_comb;
  assign p1_or_11451_comb = p1_shrl_11380_comb | p1_shll_11381_comb;
  assign p1_or_11452_comb = p1_shll_11382_comb | p1_shrl_11383_comb;
  assign p1_or_11453_comb = p1_shrl_11384_comb | p1_shll_11385_comb;
  assign p1_nor_11454_comb = ~(p1_not_11386_comb | p0_rs2);
  assign p1_nand_11455_comb = ~(p1_not_11386_comb & p0_rs2);
  assign p1_not_11456_comb = ~p1_xor_11387_comb;
  assign p1_xor_11457_comb = p1_rotation_1__1_comb ^ p1_rotation_2__1_comb ^ p1_shift_1_comb ^ p1_combined_1_comb ^ p1_combined_2_comb;
  assign p1_result__43_comb = p1_bit_slice_11391_comb ^ p1_bit_slice_11392_comb ^ p1_rotation_3__9_comb;
  assign p1_xor_11459_comb = p1_rotation_1__2_comb ^ p1_rotation_2__2_comb ^ p1_rotation_3__1_comb ^ p1_combined_1__1_comb ^ p1_combined_2__1_comb ^ p1_rotation_3__1_comb ^ p0_rs2;
  assign p1_result__23_comb = p0_rs1[25];
  assign p1_result__25_comb = p0_rs1[26];
  assign p1_result__27_comb = p0_rs1[27];
  assign p1_result__29_comb = p0_rs1[28];
  assign p1_result__31_comb = p0_rs1[29];
  assign p1_result__33_comb = p0_rs1[30];
  assign p1_result__35_comb = p0_rs1[31];
  assign p1_result__34_comb = p0_rs1[15];
  assign p1_result__32_comb = p0_rs1[14];
  assign p1_result__30_comb = p0_rs1[13];
  assign p1_result__28_comb = p0_rs1[12];
  assign p1_result__19_comb = p0_rs1[23];
  assign p1_result__15_comb = p0_rs1[21];
  assign p1_result__11_comb = p0_rs1[19];
  assign p1_result__7_comb = p0_rs1[17];
  assign p1_bit_slice_11475_comb = p1_result__39_comb[0];
  assign p1_result__38_comb = p1_bit_slice_11398_comb ^ p1_bit_slice_11318_comb ^ p1_bit_slice_11319_comb;
  assign p1_bit_slice_11477_comb = p1_result__37_comb[20];
  assign p1_bit_slice_11478_comb = p1_xor_11400_comb[0];
  assign p1_bit_slice_11479_comb = p1_xor_11401_comb[10:5];
  assign p1_bit_slice_11480_comb = p1_xor_11402_comb[1:0];
  assign p1_xor_11481_comb = p1_bit_slice_11337_comb ^ p1_bit_slice_11403_comb ^ p1_rotation_1__11_comb;
  assign p1_bit_slice_11482_comb = p1_xor_11404_comb[10];
  assign p1_bit_slice_11483_comb = p1_xor_11405_comb[4:0];
  assign p1_bit_slice_11484_comb = p1_xor_11406_comb[4:3];
  assign p1_bit_slice_11485_comb = p1_result__47_comb[4:0];
  assign p1_bit_slice_11486_comb = p1_result__46_comb[9:8];
  assign p1_bit_slice_11487_comb = p1_xor_11409_comb[4:0];
  assign p1_bit_slice_11488_comb = p1_xor_11410_comb[12:11];
  assign p1_or_11489_comb = p1_eq_11411_comb | p1_eq_11372_comb;
  assign p1_result__9_comb = p0_rs1[18];
  assign p1_result__13_comb = p0_rs1[20];
  assign p1_result__17_comb = p0_rs1[22];
  assign p1_result__26_comb = p0_rs1[11];
  assign p1_result__24_comb = p0_rs1[10];
  assign p1_result__22_comb = p0_rs1[9];
  assign p1_result__21_comb = p0_rs1[24];
  assign p1_result__18_comb = p0_rs1[7];
  assign p1_result__14_comb = p0_rs1[5];
  assign p1_result__10_comb = p0_rs1[3];
  assign p1_bit_slice_11500_comb = p1_xor_11401_comb[3:0];
  assign p1_bit_slice_11501_comb = p1_xor_11412_comb[8:7];
  assign p1_bit_slice_11502_comb = p1_xor_11406_comb[1:0];
  assign p1_bit_slice_11503_comb = p1_xor_11413_comb[13:10];
  assign p1_result__42_comb = p1_bit_slice_11319_comb ^ p1_bit_slice_11414_comb ^ p1_bit_slice_11415_comb;
  assign p1_bit_slice_11505_comb = p1_result__41_comb[3];
  assign p1_bit_slice_11506_comb = p1_xor_11417_comb[0];
  assign p1_bit_slice_11507_comb = p1_xor_11418_comb[6:2];
  assign p1_or_11508_comb = p1_eq_11411_comb | p1_eq_11371_comb;
  assign p1_bit_slice_11509_comb = p0_rs2[0];
  assign p1_literal_11510_comb = 1'h0;
  assign p1_bit_slice_11511_comb = p0_rs2[7];
  assign p1_result__20_comb = p0_rs1[8];
  assign p1_result__6_comb = p0_rs1[1];
  assign p1_bit_slice_11514_comb = p1_result__46_comb[0];
  assign p1_bit_slice_11515_comb = p1_result__45_comb[6];
  assign p1_result__16_comb = p0_rs1[6];
  assign p1_bit_slice_11517_comb = p1_xor_11412_comb[4:0];
  assign p1_bit_slice_11518_comb = p1_xor_11420_comb[9];
  assign p1_bit_slice_11519_comb = p1_xor_11404_comb[0];
  assign p1_bit_slice_11520_comb = p1_xor_11421_comb[13:9];
  assign p1_bit_slice_11521_comb = p1_result__41_comb[0];
  assign p1_bit_slice_11522_comb = p1_result__40_comb[13:9];
  assign p1_bit_slice_11523_comb = p1_xor_11410_comb[1:0];
  assign p1_bit_slice_11524_comb = p1_xor_11423_comb[9:6];
  assign p1_xor_11525_comb = p1_bit_slice_11424_comb ^ p1_rotation_2__12_comb ^ p1_bit_slice_11425_comb;
  assign p1_bit_slice_11526_comb = p1_xor_11426_comb[12:9];
  assign p1_result__44_comb = p1_bit_slice_11427_comb ^ p1_bit_slice_11428_comb ^ p1_bit_slice_11332_comb;
  assign p1_result__8_comb = p0_rs1[2];
  assign p1_result__12_comb = p0_rs1[4];
  assign p1_result__5_comb = p0_rs1[16];
  assign p1_bit_slice_11531_comb = p1_result__37_comb[3:0];
  assign p1_bit_slice_11532_comb = p1_result__36_comb[3:1];
  assign p1_bit_slice_11533_comb = p1_xor_11413_comb[0];
  assign p1_bit_slice_11534_comb = p1_xor_11430_comb[6:1];
  assign p1_bit_slice_11535_comb = p1_xor_11423_comb[4:0];
  assign p1_bit_slice_11536_comb = p1_xor_11431_comb[2:1];
  assign p1_or_11537_comb = p1_or_11432_comb | p1_eq_11371_comb | p1_eq_11372_comb;
  assign p1_concat_11538_comb = {p1_eq_11433_comb, p1_eq_11434_comb, p1_eq_11435_comb, p1_eq_11436_comb, p1_eq_11437_comb, p1_eq_11438_comb, p1_eq_11439_comb, p1_eq_11440_comb, p1_eq_11441_comb, p1_eq_11442_comb, p1_or_11443_comb, p1_eq_11411_comb, p1_eq_11444_comb, p1_eq_11359_comb, p1_eq_11445_comb, p1_eq_11446_comb, p1_eq_11447_comb, p1_eq_11448_comb, p1_eq_11449_comb, p1_eq_11450_comb};
  assign p1_bit_slice_11539_comb = p1_or_11451_comb[31];
  assign p1_bit_slice_11540_comb = p1_or_11452_comb[31];
  assign p1_bit_slice_11541_comb = p1_or_11453_comb[31];
  assign p1_bit_slice_11542_comb = p1_nor_11454_comb[31];
  assign p1_bit_slice_11543_comb = p1_nand_11455_comb[31];
  assign p1_bit_slice_11544_comb = p1_not_11456_comb[31];
  assign p1_bit_slice_11545_comb = p0_rs2[15];
  assign p1_bit_slice_11546_comb = p1_result__39_comb[1];
  assign p1_bit_slice_11547_comb = p1_xor_11400_comb[1];
  assign p1_bit_slice_11548_comb = p1_xor_11457_comb[31];
  assign p1_bit_slice_11549_comb = p1_xor_11402_comb[2];
  assign p1_bit_slice_11550_comb = p1_xor_11405_comb[5];
  assign p1_bit_slice_11551_comb = p1_result__43_comb[8];
  assign p1_bit_slice_11552_comb = p1_xor_11459_comb[31];
  assign p1_bit_slice_11553_comb = p1_result__47_comb[5];
  assign p1_bit_slice_11554_comb = p1_xor_11409_comb[5];
  assign p1_bit_slice_11555_comb = p1_xor_11417_comb[9];
  assign p1_concat_11556_comb = {p1_eq_11433_comb, p1_eq_11434_comb, p1_eq_11435_comb, p1_eq_11436_comb, p1_eq_11437_comb, p1_eq_11438_comb, p1_eq_11439_comb, p1_eq_11440_comb, p1_eq_11441_comb, p1_eq_11442_comb, p1_eq_11372_comb, p1_eq_11371_comb, p1_eq_11411_comb, p1_eq_11444_comb, p1_eq_11359_comb, p1_eq_11445_comb, p1_eq_11446_comb, p1_eq_11447_comb, p1_eq_11448_comb, p1_eq_11449_comb, p1_eq_11450_comb};
  assign p1_bit_slice_11557_comb = p1_or_11451_comb[30:24];
  assign p1_bit_slice_11558_comb = p1_or_11452_comb[30:24];
  assign p1_bit_slice_11559_comb = p1_or_11453_comb[30:24];
  assign p1_bit_slice_11560_comb = p1_nor_11454_comb[30:24];
  assign p1_bit_slice_11561_comb = p1_nand_11455_comb[30:24];
  assign p1_bit_slice_11562_comb = p1_not_11456_comb[30:24];
  assign p1_bit_slice_11563_comb = p0_rs2[14:8];
  assign p1_concat_11564_comb = {p1_result__23_comb, p1_result__25_comb, p1_result__27_comb, p1_result__29_comb, p1_result__31_comb, p1_result__33_comb, p1_result__35_comb};
  assign p1_concat_11565_comb = {p1_result__34_comb, p1_result__33_comb, p1_result__32_comb, p1_result__31_comb, p1_result__30_comb, p1_result__29_comb, p1_result__28_comb};
  assign p1_concat_11566_comb = {p1_result__31_comb, p1_result__27_comb, p1_result__23_comb, p1_result__19_comb, p1_result__15_comb, p1_result__11_comb, p1_result__7_comb};
  assign p1_concat_11567_comb = {p1_bit_slice_11475_comb, p1_result__38_comb, p1_bit_slice_11477_comb};
  assign p1_concat_11568_comb = {p1_bit_slice_11478_comb, p1_bit_slice_11479_comb};
  assign p1_bit_slice_11569_comb = p1_xor_11457_comb[30:24];
  assign p1_concat_11570_comb = {p1_bit_slice_11480_comb, p1_xor_11481_comb, p1_bit_slice_11482_comb};
  assign p1_concat_11571_comb = {p1_bit_slice_11483_comb, p1_bit_slice_11484_comb};
  assign p1_bit_slice_11572_comb = p1_result__43_comb[7:1];
  assign p1_bit_slice_11573_comb = p1_xor_11459_comb[30:24];
  assign p1_concat_11574_comb = {p1_bit_slice_11485_comb, p1_bit_slice_11486_comb};
  assign p1_concat_11575_comb = {p1_bit_slice_11487_comb, p1_bit_slice_11488_comb};
  assign p1_bit_slice_11576_comb = p1_xor_11417_comb[8:2];
  assign p1_concat_11577_comb = {p1_eq_11433_comb, p1_eq_11434_comb, p1_eq_11435_comb, p1_eq_11436_comb, p1_eq_11437_comb, p1_eq_11438_comb, p1_eq_11439_comb, p1_eq_11440_comb, p1_eq_11441_comb, p1_eq_11442_comb, p1_eq_11371_comb, p1_or_11489_comb, p1_eq_11444_comb, p1_eq_11359_comb, p1_eq_11445_comb, p1_eq_11446_comb, p1_eq_11447_comb, p1_eq_11448_comb, p1_eq_11449_comb, p1_eq_11450_comb};
  assign p1_bit_slice_11578_comb = p1_or_11451_comb[23];
  assign p1_bit_slice_11579_comb = p1_or_11452_comb[23];
  assign p1_bit_slice_11580_comb = p1_or_11453_comb[23];
  assign p1_bit_slice_11581_comb = p1_nor_11454_comb[23];
  assign p1_bit_slice_11582_comb = p1_nand_11455_comb[23];
  assign p1_bit_slice_11583_comb = p1_not_11456_comb[23];
  assign p1_bit_slice_11584_comb = p1_result__37_comb[19];
  assign p1_bit_slice_11585_comb = p1_xor_11401_comb[4];
  assign p1_bit_slice_11586_comb = p1_xor_11457_comb[23];
  assign p1_bit_slice_11587_comb = p1_xor_11404_comb[9];
  assign p1_bit_slice_11588_comb = p1_xor_11406_comb[2];
  assign p1_bit_slice_11589_comb = p1_result__43_comb[0];
  assign p1_bit_slice_11590_comb = p1_xor_11459_comb[23];
  assign p1_bit_slice_11591_comb = p1_result__46_comb[7];
  assign p1_bit_slice_11592_comb = p1_xor_11410_comb[10];
  assign p1_bit_slice_11593_comb = p1_xor_11417_comb[1];
  assign p1_bit_slice_11594_comb = p1_or_11451_comb[22:17];
  assign p1_bit_slice_11595_comb = p1_or_11452_comb[22:17];
  assign p1_bit_slice_11596_comb = p1_or_11453_comb[22:17];
  assign p1_bit_slice_11597_comb = p1_nor_11454_comb[22:17];
  assign p1_bit_slice_11598_comb = p1_nand_11455_comb[22:17];
  assign p1_bit_slice_11599_comb = p1_not_11456_comb[22:17];
  assign p1_bit_slice_11600_comb = p0_rs2[6:1];
  assign p1_concat_11601_comb = {p1_result__7_comb, p1_result__9_comb, p1_result__11_comb, p1_result__13_comb, p1_result__15_comb, p1_result__17_comb};
  assign p1_bit_slice_11602_comb = p0_rs1[14:9];
  assign p1_concat_11603_comb = {p1_result__26_comb, p1_result__25_comb, p1_result__24_comb, p1_result__23_comb, p1_result__22_comb, p1_result__21_comb};
  assign p1_concat_11604_comb = {p1_result__30_comb, p1_result__26_comb, p1_result__22_comb, p1_result__18_comb, p1_result__14_comb, p1_result__10_comb};
  assign p1_bit_slice_11605_comb = p1_result__37_comb[18:13];
  assign p1_concat_11606_comb = {p1_bit_slice_11500_comb, p1_bit_slice_11501_comb};
  assign p1_bit_slice_11607_comb = p1_xor_11457_comb[22:17];
  assign p1_bit_slice_11608_comb = p1_xor_11404_comb[8:3];
  assign p1_concat_11609_comb = {p1_bit_slice_11502_comb, p1_bit_slice_11503_comb};
  assign p1_concat_11610_comb = {p1_result__42_comb, p1_bit_slice_11505_comb};
  assign p1_bit_slice_11611_comb = p1_xor_11459_comb[22:17];
  assign p1_bit_slice_11612_comb = p1_result__46_comb[6:1];
  assign p1_bit_slice_11613_comb = p1_xor_11410_comb[9:4];
  assign p1_concat_11614_comb = {p1_bit_slice_11506_comb, p1_bit_slice_11507_comb};
  assign p1_concat_11615_comb = {p1_eq_11433_comb, p1_eq_11434_comb, p1_eq_11435_comb, p1_eq_11436_comb, p1_eq_11437_comb, p1_eq_11438_comb, p1_eq_11439_comb, p1_eq_11440_comb, p1_eq_11441_comb, p1_eq_11442_comb, p1_eq_11372_comb, p1_or_11508_comb, p1_eq_11444_comb, p1_eq_11360_comb, p1_eq_11359_comb, p1_eq_11445_comb, p1_eq_11446_comb, p1_eq_11447_comb, p1_eq_11448_comb, p1_eq_11449_comb, p1_eq_11450_comb};
  assign p1_bit_slice_11616_comb = p1_or_11451_comb[16:15];
  assign p1_bit_slice_11617_comb = p1_or_11452_comb[16:15];
  assign p1_bit_slice_11618_comb = p1_or_11453_comb[16:15];
  assign p1_bit_slice_11619_comb = p1_nor_11454_comb[16:15];
  assign p1_bit_slice_11620_comb = p1_nand_11455_comb[16:15];
  assign p1_bit_slice_11621_comb = p1_not_11456_comb[16:15];
  assign p1_concat_11622_comb = {p1_bit_slice_11509_comb, p1_result__34_comb};
  assign p1_concat_11623_comb = {p1_literal_11510_comb, p1_bit_slice_11511_comb};
  assign p1_concat_11624_comb = {p1_result__19_comb, p1_result__20_comb};
  assign p1_concat_11625_comb = {p1_result__20_comb, p1_result__19_comb};
  assign p1_concat_11626_comb = {p1_result__6_comb, p1_result__33_comb};
  assign p1_bit_slice_11627_comb = p1_result__37_comb[12:11];
  assign p1_bit_slice_11628_comb = p1_xor_11412_comb[6:5];
  assign p1_bit_slice_11629_comb = p1_xor_11457_comb[16:15];
  assign p1_bit_slice_11630_comb = p1_xor_11404_comb[2:1];
  assign p1_bit_slice_11631_comb = p1_xor_11413_comb[9:8];
  assign p1_bit_slice_11632_comb = p1_result__41_comb[2:1];
  assign p1_bit_slice_11633_comb = p1_xor_11459_comb[16:15];
  assign p1_concat_11634_comb = {p1_bit_slice_11514_comb, p1_bit_slice_11515_comb};
  assign p1_bit_slice_11635_comb = p1_xor_11410_comb[3:2];
  assign p1_bit_slice_11636_comb = p1_xor_11418_comb[1:0];
  assign p1_concat_11637_comb = {p1_eq_11433_comb, p1_eq_11434_comb, p1_eq_11435_comb, p1_eq_11436_comb, p1_eq_11437_comb, p1_eq_11438_comb, p1_eq_11439_comb, p1_eq_11440_comb, p1_eq_11441_comb, p1_eq_11442_comb, p1_eq_11372_comb, p1_eq_11371_comb, p1_eq_11411_comb, p1_eq_11444_comb, p1_eq_11360_comb, p1_eq_11359_comb, p1_eq_11445_comb, p1_eq_11446_comb, p1_eq_11447_comb, p1_eq_11448_comb, p1_eq_11449_comb, p1_eq_11450_comb};
  assign p1_bit_slice_11638_comb = p1_or_11451_comb[14:9];
  assign p1_bit_slice_11639_comb = p1_or_11452_comb[14:9];
  assign p1_bit_slice_11640_comb = p1_or_11453_comb[14:9];
  assign p1_bit_slice_11641_comb = p1_nor_11454_comb[14:9];
  assign p1_bit_slice_11642_comb = p1_nand_11455_comb[14:9];
  assign p1_bit_slice_11643_comb = p1_not_11456_comb[14:9];
  assign p1_concat_11644_comb = {p1_result__22_comb, p1_result__24_comb, p1_result__26_comb, p1_result__28_comb, p1_result__30_comb, p1_result__32_comb};
  assign p1_bit_slice_11645_comb = p0_rs1[22:17];
  assign p1_concat_11646_comb = {p1_result__18_comb, p1_result__17_comb, p1_result__16_comb, p1_result__15_comb, p1_result__14_comb, p1_result__13_comb};
  assign p1_concat_11647_comb = {p1_result__29_comb, p1_result__25_comb, p1_result__21_comb, p1_result__17_comb, p1_result__13_comb, p1_result__9_comb};
  assign p1_bit_slice_11648_comb = p1_result__37_comb[10:5];
  assign p1_concat_11649_comb = {p1_bit_slice_11517_comb, p1_bit_slice_11518_comb};
  assign p1_bit_slice_11650_comb = p1_xor_11457_comb[14:9];
  assign p1_concat_11651_comb = {p1_bit_slice_11519_comb, p1_bit_slice_11520_comb};
  assign p1_bit_slice_11652_comb = p1_xor_11413_comb[7:2];
  assign p1_concat_11653_comb = {p1_bit_slice_11521_comb, p1_bit_slice_11522_comb};
  assign p1_bit_slice_11654_comb = p1_xor_11459_comb[14:9];
  assign p1_bit_slice_11655_comb = p1_result__45_comb[5:0];
  assign p1_concat_11656_comb = {p1_bit_slice_11523_comb, p1_bit_slice_11524_comb};
  assign p1_concat_11657_comb = {p1_xor_11525_comb, p1_bit_slice_11526_comb};
  assign p1_concat_11658_comb = {p1_eq_11433_comb, p1_eq_11434_comb, p1_eq_11435_comb, p1_eq_11436_comb, p1_eq_11437_comb, p1_eq_11438_comb, p1_eq_11439_comb, p1_eq_11440_comb, p1_eq_11441_comb, p1_eq_11442_comb, p1_eq_11371_comb, p1_or_11489_comb, p1_eq_11444_comb, p1_eq_11360_comb, p1_eq_11359_comb, p1_eq_11445_comb, p1_eq_11446_comb, p1_eq_11447_comb, p1_eq_11448_comb, p1_eq_11449_comb, p1_eq_11450_comb};
  assign p1_bit_slice_11659_comb = p1_or_11451_comb[8];
  assign p1_bit_slice_11660_comb = p1_or_11452_comb[8];
  assign p1_bit_slice_11661_comb = p1_or_11453_comb[8];
  assign p1_bit_slice_11662_comb = p1_nor_11454_comb[8];
  assign p1_bit_slice_11663_comb = p1_nand_11455_comb[8];
  assign p1_bit_slice_11664_comb = p1_not_11456_comb[8];
  assign p1_bit_slice_11665_comb = p1_result__37_comb[4];
  assign p1_bit_slice_11666_comb = p1_xor_11420_comb[8];
  assign p1_bit_slice_11667_comb = p1_xor_11457_comb[8];
  assign p1_bit_slice_11668_comb = p1_xor_11421_comb[8];
  assign p1_bit_slice_11669_comb = p1_xor_11413_comb[1];
  assign p1_bit_slice_11670_comb = p1_result__40_comb[8];
  assign p1_bit_slice_11671_comb = p1_xor_11459_comb[8];
  assign p1_bit_slice_11672_comb = p1_result__44_comb[8];
  assign p1_bit_slice_11673_comb = p1_xor_11423_comb[5];
  assign p1_bit_slice_11674_comb = p1_xor_11426_comb[8];
  assign p1_concat_11675_comb = {p1_eq_11433_comb, p1_eq_11434_comb, p1_eq_11435_comb, p1_eq_11436_comb, p1_eq_11437_comb, p1_eq_11438_comb, p1_eq_11439_comb, p1_eq_11440_comb, p1_eq_11441_comb, p1_eq_11442_comb, p1_eq_11372_comb, p1_eq_11371_comb, p1_eq_11411_comb, p1_eq_11444_comb, p1_or_11432_comb, p1_eq_11445_comb, p1_eq_11446_comb, p1_eq_11447_comb, p1_eq_11448_comb, p1_eq_11449_comb, p1_eq_11450_comb};
  assign p1_bit_slice_11676_comb = p1_or_11451_comb[7:1];
  assign p1_bit_slice_11677_comb = p1_or_11452_comb[7:1];
  assign p1_bit_slice_11678_comb = p1_or_11453_comb[7:1];
  assign p1_bit_slice_11679_comb = p1_nor_11454_comb[7:1];
  assign p1_bit_slice_11680_comb = p1_nand_11455_comb[7:1];
  assign p1_bit_slice_11681_comb = p1_not_11456_comb[7:1];
  assign p1_bit_slice_11682_comb = p0_rs1[7:1];
  assign p1_concat_11683_comb = {p1_rotation_1__8_comb, p1_result__6_comb, p1_result__8_comb, p1_result__10_comb, p1_result__12_comb, p1_result__14_comb, p1_result__16_comb};
  assign p1_concat_11684_comb = {p1_result__11_comb, p1_result__10_comb, p1_result__9_comb, p1_result__8_comb, p1_result__7_comb, p1_result__6_comb, p1_result__5_comb};
  assign p1_concat_11685_comb = {p1_result__32_comb, p1_result__28_comb, p1_result__24_comb, p1_result__20_comb, p1_result__16_comb, p1_result__12_comb, p1_result__8_comb};
  assign p1_concat_11686_comb = {p1_bit_slice_11531_comb, p1_bit_slice_11532_comb};
  assign p1_bit_slice_11687_comb = p1_xor_11420_comb[7:1];
  assign p1_bit_slice_11688_comb = p1_xor_11457_comb[7:1];
  assign p1_bit_slice_11689_comb = p1_xor_11421_comb[7:1];
  assign p1_concat_11690_comb = {p1_bit_slice_11533_comb, p1_bit_slice_11534_comb};
  assign p1_bit_slice_11691_comb = p1_result__40_comb[7:1];
  assign p1_bit_slice_11692_comb = p1_xor_11459_comb[7:1];
  assign p1_bit_slice_11693_comb = p1_result__44_comb[7:1];
  assign p1_concat_11694_comb = {p1_bit_slice_11535_comb, p1_bit_slice_11536_comb};
  assign p1_bit_slice_11695_comb = p1_xor_11426_comb[7:1];
  assign p1_concat_11696_comb = {p1_eq_11433_comb, p1_eq_11434_comb, p1_eq_11435_comb, p1_eq_11436_comb, p1_eq_11437_comb, p1_eq_11438_comb, p1_eq_11439_comb, p1_eq_11440_comb, p1_eq_11441_comb, p1_eq_11442_comb, p1_eq_11411_comb, p1_eq_11444_comb, p1_or_11537_comb, p1_eq_11445_comb, p1_eq_11446_comb, p1_eq_11447_comb, p1_eq_11448_comb, p1_eq_11449_comb, p1_eq_11450_comb};
  assign p1_bit_slice_11697_comb = p1_or_11451_comb[0];
  assign p1_bit_slice_11698_comb = p1_or_11452_comb[0];
  assign p1_bit_slice_11699_comb = p1_or_11453_comb[0];
  assign p1_bit_slice_11700_comb = p1_nor_11454_comb[0];
  assign p1_bit_slice_11701_comb = p1_nand_11455_comb[0];
  assign p1_bit_slice_11702_comb = p1_not_11456_comb[0];
  assign p1_bit_slice_11703_comb = p1_result__36_comb[0];
  assign p1_bit_slice_11704_comb = p1_xor_11420_comb[0];
  assign p1_bit_slice_11705_comb = p1_xor_11457_comb[0];
  assign p1_bit_slice_11706_comb = p1_xor_11421_comb[0];
  assign p1_bit_slice_11707_comb = p1_xor_11430_comb[0];
  assign p1_bit_slice_11708_comb = p1_result__40_comb[0];
  assign p1_bit_slice_11709_comb = p1_xor_11459_comb[0];
  assign p1_bit_slice_11710_comb = p1_result__44_comb[0];
  assign p1_bit_slice_11711_comb = p1_xor_11431_comb[0];
  assign p1_bit_slice_11712_comb = p1_xor_11426_comb[0];
  assign p1_one_hot_sel_11713_comb = p1_bit_slice_11539_comb & p1_concat_11538_comb[0] | p1_bit_slice_11540_comb & p1_concat_11538_comb[1] | p1_bit_slice_11541_comb & p1_concat_11538_comb[2] | p1_bit_slice_11542_comb & p1_concat_11538_comb[3] | p1_bit_slice_11543_comb & p1_concat_11538_comb[4] | p1_bit_slice_11544_comb & p1_concat_11538_comb[5] | p1_bit_slice_11545_comb & p1_concat_11538_comb[6] | p1_result__21_comb & p1_concat_11538_comb[7] | p1_result__18_comb & p1_concat_11538_comb[8] | p1_result__35_comb & p1_concat_11538_comb[9] | p1_bit_slice_11546_comb & p1_concat_11538_comb[10] | p1_bit_slice_11547_comb & p1_concat_11538_comb[11] | p1_bit_slice_11548_comb & p1_concat_11538_comb[12] | p1_bit_slice_11549_comb & p1_concat_11538_comb[13] | p1_bit_slice_11550_comb & p1_concat_11538_comb[14] | p1_bit_slice_11551_comb & p1_concat_11538_comb[15] | p1_bit_slice_11552_comb & p1_concat_11538_comb[16] | p1_bit_slice_11553_comb & p1_concat_11538_comb[17] | p1_bit_slice_11554_comb & p1_concat_11538_comb[18] | p1_bit_slice_11555_comb & p1_concat_11538_comb[19];
  assign p1_one_hot_sel_11714_comb = p1_bit_slice_11557_comb & {7{p1_concat_11556_comb[0]}} | p1_bit_slice_11558_comb & {7{p1_concat_11556_comb[1]}} | p1_bit_slice_11559_comb & {7{p1_concat_11556_comb[2]}} | p1_bit_slice_11560_comb & {7{p1_concat_11556_comb[3]}} | p1_bit_slice_11561_comb & {7{p1_concat_11556_comb[4]}} | p1_bit_slice_11562_comb & {7{p1_concat_11556_comb[5]}} | p1_bit_slice_11563_comb & {7{p1_concat_11556_comb[6]}} | p1_concat_11564_comb & {7{p1_concat_11556_comb[7]}} | p1_rotation_3__5_comb & {7{p1_concat_11556_comb[8]}} | p1_concat_11565_comb & {7{p1_concat_11556_comb[9]}} | p1_concat_11566_comb & {7{p1_concat_11556_comb[10]}} | p1_concat_11567_comb & {7{p1_concat_11556_comb[11]}} | p1_concat_11568_comb & {7{p1_concat_11556_comb[12]}} | p1_bit_slice_11569_comb & {7{p1_concat_11556_comb[13]}} | p1_concat_11570_comb & {7{p1_concat_11556_comb[14]}} | p1_concat_11571_comb & {7{p1_concat_11556_comb[15]}} | p1_bit_slice_11572_comb & {7{p1_concat_11556_comb[16]}} | p1_bit_slice_11573_comb & {7{p1_concat_11556_comb[17]}} | p1_concat_11574_comb & {7{p1_concat_11556_comb[18]}} | p1_concat_11575_comb & {7{p1_concat_11556_comb[19]}} | p1_bit_slice_11576_comb & {7{p1_concat_11556_comb[20]}};
  assign p1_one_hot_sel_11715_comb = p1_bit_slice_11578_comb & p1_concat_11577_comb[0] | p1_bit_slice_11579_comb & p1_concat_11577_comb[1] | p1_bit_slice_11580_comb & p1_concat_11577_comb[2] | p1_bit_slice_11581_comb & p1_concat_11577_comb[3] | p1_bit_slice_11582_comb & p1_concat_11577_comb[4] | p1_bit_slice_11583_comb & p1_concat_11577_comb[5] | p1_bit_slice_11511_comb & p1_concat_11577_comb[6] | p1_result__5_comb & p1_concat_11577_comb[7] | p1_result__34_comb & p1_concat_11577_comb[8] | p1_result__27_comb & p1_concat_11577_comb[9] | p1_bit_slice_11584_comb & p1_concat_11577_comb[10] | p1_bit_slice_11585_comb & p1_concat_11577_comb[11] | p1_bit_slice_11586_comb & p1_concat_11577_comb[12] | p1_bit_slice_11587_comb & p1_concat_11577_comb[13] | p1_bit_slice_11588_comb & p1_concat_11577_comb[14] | p1_bit_slice_11589_comb & p1_concat_11577_comb[15] | p1_bit_slice_11590_comb & p1_concat_11577_comb[16] | p1_bit_slice_11591_comb & p1_concat_11577_comb[17] | p1_bit_slice_11592_comb & p1_concat_11577_comb[18] | p1_bit_slice_11593_comb & p1_concat_11577_comb[19];
  assign p1_one_hot_sel_11716_comb = p1_bit_slice_11594_comb & {6{p1_concat_11556_comb[0]}} | p1_bit_slice_11595_comb & {6{p1_concat_11556_comb[1]}} | p1_bit_slice_11596_comb & {6{p1_concat_11556_comb[2]}} | p1_bit_slice_11597_comb & {6{p1_concat_11556_comb[3]}} | p1_bit_slice_11598_comb & {6{p1_concat_11556_comb[4]}} | p1_bit_slice_11599_comb & {6{p1_concat_11556_comb[5]}} | p1_bit_slice_11600_comb & {6{p1_concat_11556_comb[6]}} | p1_concat_11601_comb & {6{p1_concat_11556_comb[7]}} | p1_bit_slice_11602_comb & {6{p1_concat_11556_comb[8]}} | p1_concat_11603_comb & {6{p1_concat_11556_comb[9]}} | p1_concat_11604_comb & {6{p1_concat_11556_comb[10]}} | p1_bit_slice_11605_comb & {6{p1_concat_11556_comb[11]}} | p1_concat_11606_comb & {6{p1_concat_11556_comb[12]}} | p1_bit_slice_11607_comb & {6{p1_concat_11556_comb[13]}} | p1_bit_slice_11608_comb & {6{p1_concat_11556_comb[14]}} | p1_concat_11609_comb & {6{p1_concat_11556_comb[15]}} | p1_concat_11610_comb & {6{p1_concat_11556_comb[16]}} | p1_bit_slice_11611_comb & {6{p1_concat_11556_comb[17]}} | p1_bit_slice_11612_comb & {6{p1_concat_11556_comb[18]}} | p1_bit_slice_11613_comb & {6{p1_concat_11556_comb[19]}} | p1_concat_11614_comb & {6{p1_concat_11556_comb[20]}};
  assign p1_one_hot_sel_11717_comb = p1_bit_slice_11616_comb & {2{p1_concat_11615_comb[0]}} | p1_bit_slice_11617_comb & {2{p1_concat_11615_comb[1]}} | p1_bit_slice_11618_comb & {2{p1_concat_11615_comb[2]}} | p1_bit_slice_11619_comb & {2{p1_concat_11615_comb[3]}} | p1_bit_slice_11620_comb & {2{p1_concat_11615_comb[4]}} | p1_bit_slice_11621_comb & {2{p1_concat_11615_comb[5]}} | p1_concat_11622_comb & {2{p1_concat_11615_comb[6]}} | p1_concat_11623_comb & {2{p1_concat_11615_comb[7]}} | p1_concat_11624_comb & {2{p1_concat_11615_comb[8]}} | p1_concat_11625_comb & {2{p1_concat_11615_comb[9]}} | p1_concat_11626_comb & {2{p1_concat_11615_comb[10]}} | p1_bit_slice_11627_comb & {2{p1_concat_11615_comb[11]}} | p1_bit_slice_11628_comb & {2{p1_concat_11615_comb[12]}} | p1_bit_slice_11629_comb & {2{p1_concat_11615_comb[13]}} | p1_bit_slice_11630_comb & {2{p1_concat_11615_comb[14]}} | p1_bit_slice_11631_comb & {2{p1_concat_11615_comb[15]}} | p1_bit_slice_11632_comb & {2{p1_concat_11615_comb[16]}} | p1_bit_slice_11633_comb & {2{p1_concat_11615_comb[17]}} | p1_concat_11634_comb & {2{p1_concat_11615_comb[18]}} | p1_bit_slice_11635_comb & {2{p1_concat_11615_comb[19]}} | p1_bit_slice_11636_comb & {2{p1_concat_11615_comb[20]}};
  assign p1_one_hot_sel_11718_comb = p1_bit_slice_11638_comb & {6{p1_concat_11637_comb[0]}} | p1_bit_slice_11639_comb & {6{p1_concat_11637_comb[1]}} | p1_bit_slice_11640_comb & {6{p1_concat_11637_comb[2]}} | p1_bit_slice_11641_comb & {6{p1_concat_11637_comb[3]}} | p1_bit_slice_11642_comb & {6{p1_concat_11637_comb[4]}} | p1_bit_slice_11643_comb & {6{p1_concat_11637_comb[5]}} | p1_bit_slice_11602_comb & {6{p1_concat_11637_comb[6]}} | p1_bit_slice_11600_comb & {6{p1_concat_11637_comb[7]}} | p1_concat_11644_comb & {6{p1_concat_11637_comb[8]}} | p1_bit_slice_11645_comb & {6{p1_concat_11637_comb[9]}} | p1_concat_11646_comb & {6{p1_concat_11637_comb[10]}} | p1_concat_11647_comb & {6{p1_concat_11637_comb[11]}} | p1_bit_slice_11648_comb & {6{p1_concat_11637_comb[12]}} | p1_concat_11649_comb & {6{p1_concat_11637_comb[13]}} | p1_bit_slice_11650_comb & {6{p1_concat_11637_comb[14]}} | p1_concat_11651_comb & {6{p1_concat_11637_comb[15]}} | p1_bit_slice_11652_comb & {6{p1_concat_11637_comb[16]}} | p1_concat_11653_comb & {6{p1_concat_11637_comb[17]}} | p1_bit_slice_11654_comb & {6{p1_concat_11637_comb[18]}} | p1_bit_slice_11655_comb & {6{p1_concat_11637_comb[19]}} | p1_concat_11656_comb & {6{p1_concat_11637_comb[20]}} | p1_concat_11657_comb & {6{p1_concat_11637_comb[21]}};
  assign p1_one_hot_sel_11719_comb = p1_bit_slice_11659_comb & p1_concat_11658_comb[0] | p1_bit_slice_11660_comb & p1_concat_11658_comb[1] | p1_bit_slice_11661_comb & p1_concat_11658_comb[2] | p1_bit_slice_11662_comb & p1_concat_11658_comb[3] | p1_bit_slice_11663_comb & p1_concat_11658_comb[4] | p1_bit_slice_11664_comb & p1_concat_11658_comb[5] | p1_result__20_comb & p1_concat_11658_comb[6] | p1_bit_slice_11509_comb & p1_concat_11658_comb[7] | p1_result__34_comb & p1_concat_11658_comb[8] | p1_result__5_comb & p1_concat_11658_comb[9] | p1_result__12_comb & p1_concat_11658_comb[10] | p1_bit_slice_11665_comb & p1_concat_11658_comb[11] | p1_bit_slice_11666_comb & p1_concat_11658_comb[12] | p1_bit_slice_11667_comb & p1_concat_11658_comb[13] | p1_bit_slice_11668_comb & p1_concat_11658_comb[14] | p1_bit_slice_11669_comb & p1_concat_11658_comb[15] | p1_bit_slice_11670_comb & p1_concat_11658_comb[16] | p1_bit_slice_11671_comb & p1_concat_11658_comb[17] | p1_bit_slice_11672_comb & p1_concat_11658_comb[18] | p1_bit_slice_11673_comb & p1_concat_11658_comb[19] | p1_bit_slice_11674_comb & p1_concat_11658_comb[20];
  assign p1_one_hot_sel_11720_comb = p1_bit_slice_11676_comb & {7{p1_concat_11675_comb[0]}} | p1_bit_slice_11677_comb & {7{p1_concat_11675_comb[1]}} | p1_bit_slice_11678_comb & {7{p1_concat_11675_comb[2]}} | p1_bit_slice_11679_comb & {7{p1_concat_11675_comb[3]}} | p1_bit_slice_11680_comb & {7{p1_concat_11675_comb[4]}} | p1_bit_slice_11681_comb & {7{p1_concat_11675_comb[5]}} | p1_bit_slice_11682_comb & {7{p1_concat_11675_comb[6]}} | p1_concat_11683_comb & {7{p1_concat_11675_comb[7]}} | p1_rotation_3__6_comb & {7{p1_concat_11675_comb[8]}} | p1_concat_11684_comb & {7{p1_concat_11675_comb[9]}} | p1_concat_11685_comb & {7{p1_concat_11675_comb[10]}} | p1_concat_11686_comb & {7{p1_concat_11675_comb[11]}} | p1_bit_slice_11687_comb & {7{p1_concat_11675_comb[12]}} | p1_bit_slice_11688_comb & {7{p1_concat_11675_comb[13]}} | p1_bit_slice_11689_comb & {7{p1_concat_11675_comb[14]}} | p1_concat_11690_comb & {7{p1_concat_11675_comb[15]}} | p1_bit_slice_11691_comb & {7{p1_concat_11675_comb[16]}} | p1_bit_slice_11692_comb & {7{p1_concat_11675_comb[17]}} | p1_bit_slice_11693_comb & {7{p1_concat_11675_comb[18]}} | p1_concat_11694_comb & {7{p1_concat_11675_comb[19]}} | p1_bit_slice_11695_comb & {7{p1_concat_11675_comb[20]}};
  assign p1_one_hot_sel_11721_comb = p1_bit_slice_11697_comb & p1_concat_11696_comb[0] | p1_bit_slice_11698_comb & p1_concat_11696_comb[1] | p1_bit_slice_11699_comb & p1_concat_11696_comb[2] | p1_bit_slice_11700_comb & p1_concat_11696_comb[3] | p1_bit_slice_11701_comb & p1_concat_11696_comb[4] | p1_bit_slice_11702_comb & p1_concat_11696_comb[5] | p1_rotation_1__8_comb & p1_concat_11696_comb[6] | p1_result__18_comb & p1_concat_11696_comb[7] | p1_result__21_comb & p1_concat_11696_comb[8] | p1_bit_slice_11703_comb & p1_concat_11696_comb[9] | p1_bit_slice_11704_comb & p1_concat_11696_comb[10] | p1_bit_slice_11705_comb & p1_concat_11696_comb[11] | p1_bit_slice_11706_comb & p1_concat_11696_comb[12] | p1_bit_slice_11707_comb & p1_concat_11696_comb[13] | p1_bit_slice_11708_comb & p1_concat_11696_comb[14] | p1_bit_slice_11709_comb & p1_concat_11696_comb[15] | p1_bit_slice_11710_comb & p1_concat_11696_comb[16] | p1_bit_slice_11711_comb & p1_concat_11696_comb[17] | p1_bit_slice_11712_comb & p1_concat_11696_comb[18];
  assign p1_literal_11722_comb = 32'h0000_0016;
  assign p1_concat_11723_comb = {p1_one_hot_sel_11713_comb, p1_one_hot_sel_11714_comb, p1_one_hot_sel_11715_comb, p1_one_hot_sel_11716_comb, p1_one_hot_sel_11717_comb, p1_one_hot_sel_11718_comb, p1_one_hot_sel_11719_comb, p1_one_hot_sel_11720_comb, p1_one_hot_sel_11721_comb};
  assign p1_ult_11724_comb = p0_instruction < p1_literal_11722_comb;
  assign p1_tuple_11725_comb = {p1_concat_11723_comb, p1_ult_11724_comb};

  // Registers for pipe stage 1:
  reg [32:0] p1_tuple_11725;
  always_ff @ (posedge clk) begin
    p1_tuple_11725 <= p1_tuple_11725_comb;
  end
  assign out = p1_tuple_11725;
endmodule
