VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_proj_example
  CLASS BLOCK ;
  FOREIGN user_proj_example ;
  ORIGIN 0.000 0.000 ;
  SIZE 2800.000 BY 1760.000 ;
  PIN la_data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 56.210 0.000 56.490 4.000 ;
    END
  END la_data_in[0]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 479.410 0.000 479.690 4.000 ;
    END
  END la_data_in[10]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 521.730 0.000 522.010 4.000 ;
    END
  END la_data_in[11]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 564.050 0.000 564.330 4.000 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 606.370 0.000 606.650 4.000 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 648.690 0.000 648.970 4.000 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 691.010 0.000 691.290 4.000 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 733.330 0.000 733.610 4.000 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 775.650 0.000 775.930 4.000 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 817.970 0.000 818.250 4.000 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 860.290 0.000 860.570 4.000 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 98.530 0.000 98.810 4.000 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 902.610 0.000 902.890 4.000 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 944.930 0.000 945.210 4.000 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 987.250 0.000 987.530 4.000 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1029.570 0.000 1029.850 4.000 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1071.890 0.000 1072.170 4.000 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1114.210 0.000 1114.490 4.000 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1156.530 0.000 1156.810 4.000 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1198.850 0.000 1199.130 4.000 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1241.170 0.000 1241.450 4.000 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1283.490 0.000 1283.770 4.000 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 140.850 0.000 141.130 4.000 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1325.810 0.000 1326.090 4.000 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1368.130 0.000 1368.410 4.000 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1410.450 0.000 1410.730 4.000 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1452.770 0.000 1453.050 4.000 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1473.930 0.000 1474.210 4.000 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1495.090 0.000 1495.370 4.000 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1516.250 0.000 1516.530 4.000 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1537.410 0.000 1537.690 4.000 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1558.570 0.000 1558.850 4.000 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1579.730 0.000 1580.010 4.000 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 183.170 0.000 183.450 4.000 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1600.890 0.000 1601.170 4.000 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1622.050 0.000 1622.330 4.000 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1643.210 0.000 1643.490 4.000 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1664.370 0.000 1664.650 4.000 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1685.530 0.000 1685.810 4.000 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1706.690 0.000 1706.970 4.000 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1727.850 0.000 1728.130 4.000 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1749.010 0.000 1749.290 4.000 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1770.170 0.000 1770.450 4.000 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1791.330 0.000 1791.610 4.000 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 225.490 0.000 225.770 4.000 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1812.490 0.000 1812.770 4.000 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1833.650 0.000 1833.930 4.000 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1854.810 0.000 1855.090 4.000 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1875.970 0.000 1876.250 4.000 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1897.130 0.000 1897.410 4.000 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1918.290 0.000 1918.570 4.000 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1939.450 0.000 1939.730 4.000 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1960.610 0.000 1960.890 4.000 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 1981.770 0.000 1982.050 4.000 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 2002.930 0.000 2003.210 4.000 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 267.810 0.000 268.090 4.000 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 2024.090 0.000 2024.370 4.000 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 2045.250 0.000 2045.530 4.000 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 2066.410 0.000 2066.690 4.000 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 2087.570 0.000 2087.850 4.000 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 2108.730 0.000 2109.010 4.000 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 2129.890 0.000 2130.170 4.000 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 2151.050 0.000 2151.330 4.000 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 2172.210 0.000 2172.490 4.000 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 2193.370 0.000 2193.650 4.000 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 2214.530 0.000 2214.810 4.000 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 310.130 0.000 310.410 4.000 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 2235.690 0.000 2235.970 4.000 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 2256.850 0.000 2257.130 4.000 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 2278.010 0.000 2278.290 4.000 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 2299.170 0.000 2299.450 4.000 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 2320.330 0.000 2320.610 4.000 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 2341.490 0.000 2341.770 4.000 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 2362.650 0.000 2362.930 4.000 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 2383.810 0.000 2384.090 4.000 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 2404.970 0.000 2405.250 4.000 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 2426.130 0.000 2426.410 4.000 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 352.450 0.000 352.730 4.000 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 2447.290 0.000 2447.570 4.000 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 2468.450 0.000 2468.730 4.000 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 2489.610 0.000 2489.890 4.000 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 2510.770 0.000 2511.050 4.000 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 2531.930 0.000 2532.210 4.000 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 2553.090 0.000 2553.370 4.000 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 2574.250 0.000 2574.530 4.000 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 2595.410 0.000 2595.690 4.000 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 2616.570 0.000 2616.850 4.000 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 2637.730 0.000 2638.010 4.000 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 394.770 0.000 395.050 4.000 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 2658.890 0.000 2659.170 4.000 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 2680.050 0.000 2680.330 4.000 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 2701.210 0.000 2701.490 4.000 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 2722.370 0.000 2722.650 4.000 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 2743.530 0.000 2743.810 4.000 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 2764.690 0.000 2764.970 4.000 ;
    END
  END la_data_in[95]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 437.090 0.000 437.370 4.000 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 4.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 500.570 0.000 500.850 4.000 ;
    END
  END la_data_out[10]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 542.890 0.000 543.170 4.000 ;
    END
  END la_data_out[11]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 585.210 0.000 585.490 4.000 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 627.530 0.000 627.810 4.000 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 669.850 0.000 670.130 4.000 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 712.170 0.000 712.450 4.000 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 754.490 0.000 754.770 4.000 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 796.810 0.000 797.090 4.000 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 839.130 0.000 839.410 4.000 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 881.450 0.000 881.730 4.000 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 119.690 0.000 119.970 4.000 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 923.770 0.000 924.050 4.000 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 966.090 0.000 966.370 4.000 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1008.410 0.000 1008.690 4.000 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1050.730 0.000 1051.010 4.000 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1093.050 0.000 1093.330 4.000 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1135.370 0.000 1135.650 4.000 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1177.690 0.000 1177.970 4.000 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1220.010 0.000 1220.290 4.000 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1262.330 0.000 1262.610 4.000 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1304.650 0.000 1304.930 4.000 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 162.010 0.000 162.290 4.000 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1346.970 0.000 1347.250 4.000 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1389.290 0.000 1389.570 4.000 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 1431.610 0.000 1431.890 4.000 ;
    END
  END la_data_out[32]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 204.330 0.000 204.610 4.000 ;
    END
  END la_data_out[3]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 246.650 0.000 246.930 4.000 ;
    END
  END la_data_out[4]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 288.970 0.000 289.250 4.000 ;
    END
  END la_data_out[5]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 331.290 0.000 331.570 4.000 ;
    END
  END la_data_out[6]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 373.610 0.000 373.890 4.000 ;
    END
  END la_data_out[7]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 415.930 0.000 416.210 4.000 ;
    END
  END la_data_out[8]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 2.673000 ;
    PORT
      LAYER met2 ;
        RECT 458.250 0.000 458.530 4.000 ;
    END
  END la_data_out[9]
  PIN vccd1
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 942.640 10.640 944.240 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1096.240 10.640 1097.840 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1249.840 10.640 1251.440 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1403.440 10.640 1405.040 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1557.040 10.640 1558.640 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1710.640 10.640 1712.240 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1864.240 10.640 1865.840 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2017.840 10.640 2019.440 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2171.440 10.640 2173.040 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2325.040 10.640 2326.640 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2478.640 10.640 2480.240 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2632.240 10.640 2633.840 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2785.840 10.640 2787.440 1749.200 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 865.840 10.640 867.440 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1019.440 10.640 1021.040 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1173.040 10.640 1174.640 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1326.640 10.640 1328.240 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1480.240 10.640 1481.840 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1633.840 10.640 1635.440 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1787.440 10.640 1789.040 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 1941.040 10.640 1942.640 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2094.640 10.640 2096.240 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2248.240 10.640 2249.840 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2401.840 10.640 2403.440 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2555.440 10.640 2557.040 1749.200 ;
    END
    PORT
      LAYER met4 ;
        RECT 2709.040 10.640 2710.640 1749.200 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met2 ;
        RECT 35.050 0.000 35.330 4.000 ;
    END
  END wb_clk_i
  OBS
      LAYER nwell ;
        RECT 5.330 1747.545 2794.230 1749.150 ;
        RECT 5.330 1742.105 2794.230 1744.935 ;
        RECT 5.330 1736.665 2794.230 1739.495 ;
        RECT 5.330 1731.225 2794.230 1734.055 ;
        RECT 5.330 1725.785 2794.230 1728.615 ;
        RECT 5.330 1720.345 2794.230 1723.175 ;
        RECT 5.330 1714.905 2794.230 1717.735 ;
        RECT 5.330 1709.465 2794.230 1712.295 ;
        RECT 5.330 1704.025 2794.230 1706.855 ;
        RECT 5.330 1698.585 2794.230 1701.415 ;
        RECT 5.330 1693.145 2794.230 1695.975 ;
        RECT 5.330 1687.705 2794.230 1690.535 ;
        RECT 5.330 1682.265 2794.230 1685.095 ;
        RECT 5.330 1676.825 2794.230 1679.655 ;
        RECT 5.330 1671.385 2794.230 1674.215 ;
        RECT 5.330 1665.945 2794.230 1668.775 ;
        RECT 5.330 1660.505 2794.230 1663.335 ;
        RECT 5.330 1655.065 2794.230 1657.895 ;
        RECT 5.330 1649.625 2794.230 1652.455 ;
        RECT 5.330 1644.185 2794.230 1647.015 ;
        RECT 5.330 1638.745 2794.230 1641.575 ;
        RECT 5.330 1633.305 2794.230 1636.135 ;
        RECT 5.330 1627.865 2794.230 1630.695 ;
        RECT 5.330 1622.425 2794.230 1625.255 ;
        RECT 5.330 1616.985 2794.230 1619.815 ;
        RECT 5.330 1611.545 2794.230 1614.375 ;
        RECT 5.330 1606.105 2794.230 1608.935 ;
        RECT 5.330 1600.665 2794.230 1603.495 ;
        RECT 5.330 1595.225 2794.230 1598.055 ;
        RECT 5.330 1589.785 2794.230 1592.615 ;
        RECT 5.330 1584.345 2794.230 1587.175 ;
        RECT 5.330 1578.905 2794.230 1581.735 ;
        RECT 5.330 1573.465 2794.230 1576.295 ;
        RECT 5.330 1568.025 2794.230 1570.855 ;
        RECT 5.330 1562.585 2794.230 1565.415 ;
        RECT 5.330 1557.145 2794.230 1559.975 ;
        RECT 5.330 1551.705 2794.230 1554.535 ;
        RECT 5.330 1546.265 2794.230 1549.095 ;
        RECT 5.330 1540.825 2794.230 1543.655 ;
        RECT 5.330 1535.385 2794.230 1538.215 ;
        RECT 5.330 1529.945 2794.230 1532.775 ;
        RECT 5.330 1524.505 2794.230 1527.335 ;
        RECT 5.330 1519.065 2794.230 1521.895 ;
        RECT 5.330 1513.625 2794.230 1516.455 ;
        RECT 5.330 1508.185 2794.230 1511.015 ;
        RECT 5.330 1502.745 2794.230 1505.575 ;
        RECT 5.330 1497.305 2794.230 1500.135 ;
        RECT 5.330 1491.865 2794.230 1494.695 ;
        RECT 5.330 1486.425 2794.230 1489.255 ;
        RECT 5.330 1480.985 2794.230 1483.815 ;
        RECT 5.330 1475.545 2794.230 1478.375 ;
        RECT 5.330 1470.105 2794.230 1472.935 ;
        RECT 5.330 1464.665 2794.230 1467.495 ;
        RECT 5.330 1459.225 2794.230 1462.055 ;
        RECT 5.330 1453.785 2794.230 1456.615 ;
        RECT 5.330 1448.345 2794.230 1451.175 ;
        RECT 5.330 1442.905 2794.230 1445.735 ;
        RECT 5.330 1437.465 2794.230 1440.295 ;
        RECT 5.330 1432.025 2794.230 1434.855 ;
        RECT 5.330 1426.585 2794.230 1429.415 ;
        RECT 5.330 1421.145 2794.230 1423.975 ;
        RECT 5.330 1415.705 2794.230 1418.535 ;
        RECT 5.330 1410.265 2794.230 1413.095 ;
        RECT 5.330 1404.825 2794.230 1407.655 ;
        RECT 5.330 1399.385 2794.230 1402.215 ;
        RECT 5.330 1393.945 2794.230 1396.775 ;
        RECT 5.330 1388.505 2794.230 1391.335 ;
        RECT 5.330 1383.065 2794.230 1385.895 ;
        RECT 5.330 1377.625 2794.230 1380.455 ;
        RECT 5.330 1372.185 2794.230 1375.015 ;
        RECT 5.330 1366.745 2794.230 1369.575 ;
        RECT 5.330 1361.305 2794.230 1364.135 ;
        RECT 5.330 1355.865 2794.230 1358.695 ;
        RECT 5.330 1350.425 2794.230 1353.255 ;
        RECT 5.330 1344.985 2794.230 1347.815 ;
        RECT 5.330 1339.545 2794.230 1342.375 ;
        RECT 5.330 1334.105 2794.230 1336.935 ;
        RECT 5.330 1328.665 2794.230 1331.495 ;
        RECT 5.330 1323.225 2794.230 1326.055 ;
        RECT 5.330 1317.785 2794.230 1320.615 ;
        RECT 5.330 1312.345 2794.230 1315.175 ;
        RECT 5.330 1306.905 2794.230 1309.735 ;
        RECT 5.330 1301.465 2794.230 1304.295 ;
        RECT 5.330 1296.025 2794.230 1298.855 ;
        RECT 5.330 1290.585 2794.230 1293.415 ;
        RECT 5.330 1285.145 2794.230 1287.975 ;
        RECT 5.330 1279.705 2794.230 1282.535 ;
        RECT 5.330 1274.265 2794.230 1277.095 ;
        RECT 5.330 1268.825 2794.230 1271.655 ;
        RECT 5.330 1263.385 2794.230 1266.215 ;
        RECT 5.330 1257.945 2794.230 1260.775 ;
        RECT 5.330 1252.505 2794.230 1255.335 ;
        RECT 5.330 1247.065 2794.230 1249.895 ;
        RECT 5.330 1241.625 2794.230 1244.455 ;
        RECT 5.330 1236.185 2794.230 1239.015 ;
        RECT 5.330 1230.745 2794.230 1233.575 ;
        RECT 5.330 1225.305 2794.230 1228.135 ;
        RECT 5.330 1219.865 2794.230 1222.695 ;
        RECT 5.330 1214.425 2794.230 1217.255 ;
        RECT 5.330 1208.985 2794.230 1211.815 ;
        RECT 5.330 1203.545 2794.230 1206.375 ;
        RECT 5.330 1198.105 2794.230 1200.935 ;
        RECT 5.330 1192.665 2794.230 1195.495 ;
        RECT 5.330 1187.225 2794.230 1190.055 ;
        RECT 5.330 1181.785 2794.230 1184.615 ;
        RECT 5.330 1176.345 2794.230 1179.175 ;
        RECT 5.330 1170.905 2794.230 1173.735 ;
        RECT 5.330 1165.465 2794.230 1168.295 ;
        RECT 5.330 1160.025 2794.230 1162.855 ;
        RECT 5.330 1154.585 2794.230 1157.415 ;
        RECT 5.330 1149.145 2794.230 1151.975 ;
        RECT 5.330 1143.705 2794.230 1146.535 ;
        RECT 5.330 1138.265 2794.230 1141.095 ;
        RECT 5.330 1132.825 2794.230 1135.655 ;
        RECT 5.330 1127.385 2794.230 1130.215 ;
        RECT 5.330 1121.945 2794.230 1124.775 ;
        RECT 5.330 1116.505 2794.230 1119.335 ;
        RECT 5.330 1111.065 2794.230 1113.895 ;
        RECT 5.330 1105.625 2794.230 1108.455 ;
        RECT 5.330 1100.185 2794.230 1103.015 ;
        RECT 5.330 1094.745 2794.230 1097.575 ;
        RECT 5.330 1089.305 2794.230 1092.135 ;
        RECT 5.330 1083.865 2794.230 1086.695 ;
        RECT 5.330 1078.425 2794.230 1081.255 ;
        RECT 5.330 1072.985 2794.230 1075.815 ;
        RECT 5.330 1067.545 2794.230 1070.375 ;
        RECT 5.330 1062.105 2794.230 1064.935 ;
        RECT 5.330 1056.665 2794.230 1059.495 ;
        RECT 5.330 1051.225 2794.230 1054.055 ;
        RECT 5.330 1045.785 2794.230 1048.615 ;
        RECT 5.330 1040.345 2794.230 1043.175 ;
        RECT 5.330 1034.905 2794.230 1037.735 ;
        RECT 5.330 1029.465 2794.230 1032.295 ;
        RECT 5.330 1024.025 2794.230 1026.855 ;
        RECT 5.330 1018.585 2794.230 1021.415 ;
        RECT 5.330 1013.145 2794.230 1015.975 ;
        RECT 5.330 1007.705 2794.230 1010.535 ;
        RECT 5.330 1002.265 2794.230 1005.095 ;
        RECT 5.330 996.825 2794.230 999.655 ;
        RECT 5.330 991.385 2794.230 994.215 ;
        RECT 5.330 985.945 2794.230 988.775 ;
        RECT 5.330 980.505 2794.230 983.335 ;
        RECT 5.330 975.065 2794.230 977.895 ;
        RECT 5.330 969.625 2794.230 972.455 ;
        RECT 5.330 964.185 2794.230 967.015 ;
        RECT 5.330 958.745 2794.230 961.575 ;
        RECT 5.330 953.305 2794.230 956.135 ;
        RECT 5.330 947.865 2794.230 950.695 ;
        RECT 5.330 942.425 2794.230 945.255 ;
        RECT 5.330 936.985 2794.230 939.815 ;
        RECT 5.330 931.545 2794.230 934.375 ;
        RECT 5.330 926.105 2794.230 928.935 ;
        RECT 5.330 920.665 2794.230 923.495 ;
        RECT 5.330 915.225 2794.230 918.055 ;
        RECT 5.330 909.785 2794.230 912.615 ;
        RECT 5.330 904.345 2794.230 907.175 ;
        RECT 5.330 898.905 2794.230 901.735 ;
        RECT 5.330 893.465 2794.230 896.295 ;
        RECT 5.330 888.025 2794.230 890.855 ;
        RECT 5.330 882.585 2794.230 885.415 ;
        RECT 5.330 877.145 2794.230 879.975 ;
        RECT 5.330 871.705 2794.230 874.535 ;
        RECT 5.330 866.265 2794.230 869.095 ;
        RECT 5.330 860.825 2794.230 863.655 ;
        RECT 5.330 855.385 2794.230 858.215 ;
        RECT 5.330 849.945 2794.230 852.775 ;
        RECT 5.330 844.505 2794.230 847.335 ;
        RECT 5.330 839.065 2794.230 841.895 ;
        RECT 5.330 833.625 2794.230 836.455 ;
        RECT 5.330 828.185 2794.230 831.015 ;
        RECT 5.330 822.745 2794.230 825.575 ;
        RECT 5.330 817.305 2794.230 820.135 ;
        RECT 5.330 811.865 2794.230 814.695 ;
        RECT 5.330 806.425 2794.230 809.255 ;
        RECT 5.330 800.985 2794.230 803.815 ;
        RECT 5.330 795.545 2794.230 798.375 ;
        RECT 5.330 790.105 2794.230 792.935 ;
        RECT 5.330 784.665 2794.230 787.495 ;
        RECT 5.330 779.225 2794.230 782.055 ;
        RECT 5.330 773.785 2794.230 776.615 ;
        RECT 5.330 768.345 2794.230 771.175 ;
        RECT 5.330 762.905 2794.230 765.735 ;
        RECT 5.330 757.465 2794.230 760.295 ;
        RECT 5.330 752.025 2794.230 754.855 ;
        RECT 5.330 746.585 2794.230 749.415 ;
        RECT 5.330 741.145 2794.230 743.975 ;
        RECT 5.330 735.705 2794.230 738.535 ;
        RECT 5.330 730.265 2794.230 733.095 ;
        RECT 5.330 724.825 2794.230 727.655 ;
        RECT 5.330 719.385 2794.230 722.215 ;
        RECT 5.330 713.945 2794.230 716.775 ;
        RECT 5.330 708.505 2794.230 711.335 ;
        RECT 5.330 703.065 2794.230 705.895 ;
        RECT 5.330 697.625 2794.230 700.455 ;
        RECT 5.330 692.185 2794.230 695.015 ;
        RECT 5.330 686.745 2794.230 689.575 ;
        RECT 5.330 681.305 2794.230 684.135 ;
        RECT 5.330 675.865 2794.230 678.695 ;
        RECT 5.330 670.425 2794.230 673.255 ;
        RECT 5.330 664.985 2794.230 667.815 ;
        RECT 5.330 659.545 2794.230 662.375 ;
        RECT 5.330 654.105 2794.230 656.935 ;
        RECT 5.330 648.665 2794.230 651.495 ;
        RECT 5.330 643.225 2794.230 646.055 ;
        RECT 5.330 637.785 2794.230 640.615 ;
        RECT 5.330 632.345 2794.230 635.175 ;
        RECT 5.330 626.905 2794.230 629.735 ;
        RECT 5.330 621.465 2794.230 624.295 ;
        RECT 5.330 616.025 2794.230 618.855 ;
        RECT 5.330 610.585 2794.230 613.415 ;
        RECT 5.330 605.145 2794.230 607.975 ;
        RECT 5.330 599.705 2794.230 602.535 ;
        RECT 5.330 594.265 2794.230 597.095 ;
        RECT 5.330 588.825 2794.230 591.655 ;
        RECT 5.330 583.385 2794.230 586.215 ;
        RECT 5.330 577.945 2794.230 580.775 ;
        RECT 5.330 572.505 2794.230 575.335 ;
        RECT 5.330 567.065 2794.230 569.895 ;
        RECT 5.330 561.625 2794.230 564.455 ;
        RECT 5.330 556.185 2794.230 559.015 ;
        RECT 5.330 550.745 2794.230 553.575 ;
        RECT 5.330 545.305 2794.230 548.135 ;
        RECT 5.330 539.865 2794.230 542.695 ;
        RECT 5.330 534.425 2794.230 537.255 ;
        RECT 5.330 528.985 2794.230 531.815 ;
        RECT 5.330 523.545 2794.230 526.375 ;
        RECT 5.330 518.105 2794.230 520.935 ;
        RECT 5.330 512.665 2794.230 515.495 ;
        RECT 5.330 507.225 2794.230 510.055 ;
        RECT 5.330 501.785 2794.230 504.615 ;
        RECT 5.330 496.345 2794.230 499.175 ;
        RECT 5.330 490.905 2794.230 493.735 ;
        RECT 5.330 485.465 2794.230 488.295 ;
        RECT 5.330 480.025 2794.230 482.855 ;
        RECT 5.330 474.585 2794.230 477.415 ;
        RECT 5.330 469.145 2794.230 471.975 ;
        RECT 5.330 463.705 2794.230 466.535 ;
        RECT 5.330 458.265 2794.230 461.095 ;
        RECT 5.330 452.825 2794.230 455.655 ;
        RECT 5.330 447.385 2794.230 450.215 ;
        RECT 5.330 441.945 2794.230 444.775 ;
        RECT 5.330 436.505 2794.230 439.335 ;
        RECT 5.330 431.065 2794.230 433.895 ;
        RECT 5.330 425.625 2794.230 428.455 ;
        RECT 5.330 420.185 2794.230 423.015 ;
        RECT 5.330 414.745 2794.230 417.575 ;
        RECT 5.330 409.305 2794.230 412.135 ;
        RECT 5.330 403.865 2794.230 406.695 ;
        RECT 5.330 398.425 2794.230 401.255 ;
        RECT 5.330 392.985 2794.230 395.815 ;
        RECT 5.330 387.545 2794.230 390.375 ;
        RECT 5.330 382.105 2794.230 384.935 ;
        RECT 5.330 376.665 2794.230 379.495 ;
        RECT 5.330 371.225 2794.230 374.055 ;
        RECT 5.330 365.785 2794.230 368.615 ;
        RECT 5.330 360.345 2794.230 363.175 ;
        RECT 5.330 354.905 2794.230 357.735 ;
        RECT 5.330 349.465 2794.230 352.295 ;
        RECT 5.330 344.025 2794.230 346.855 ;
        RECT 5.330 338.585 2794.230 341.415 ;
        RECT 5.330 333.145 2794.230 335.975 ;
        RECT 5.330 327.705 2794.230 330.535 ;
        RECT 5.330 322.265 2794.230 325.095 ;
        RECT 5.330 316.825 2794.230 319.655 ;
        RECT 5.330 311.385 2794.230 314.215 ;
        RECT 5.330 305.945 2794.230 308.775 ;
        RECT 5.330 300.505 2794.230 303.335 ;
        RECT 5.330 295.065 2794.230 297.895 ;
        RECT 5.330 289.625 2794.230 292.455 ;
        RECT 5.330 284.185 2794.230 287.015 ;
        RECT 5.330 278.745 2794.230 281.575 ;
        RECT 5.330 273.305 2794.230 276.135 ;
        RECT 5.330 267.865 2794.230 270.695 ;
        RECT 5.330 262.425 2794.230 265.255 ;
        RECT 5.330 256.985 2794.230 259.815 ;
        RECT 5.330 251.545 2794.230 254.375 ;
        RECT 5.330 246.105 2794.230 248.935 ;
        RECT 5.330 240.665 2794.230 243.495 ;
        RECT 5.330 235.225 2794.230 238.055 ;
        RECT 5.330 229.785 2794.230 232.615 ;
        RECT 5.330 224.345 2794.230 227.175 ;
        RECT 5.330 218.905 2794.230 221.735 ;
        RECT 5.330 213.465 2794.230 216.295 ;
        RECT 5.330 208.025 2794.230 210.855 ;
        RECT 5.330 202.585 2794.230 205.415 ;
        RECT 5.330 197.145 2794.230 199.975 ;
        RECT 5.330 191.705 2794.230 194.535 ;
        RECT 5.330 186.265 2794.230 189.095 ;
        RECT 5.330 180.825 2794.230 183.655 ;
        RECT 5.330 175.385 2794.230 178.215 ;
        RECT 5.330 169.945 2794.230 172.775 ;
        RECT 5.330 164.505 2794.230 167.335 ;
        RECT 5.330 159.065 2794.230 161.895 ;
        RECT 5.330 153.625 2794.230 156.455 ;
        RECT 5.330 148.185 2794.230 151.015 ;
        RECT 5.330 142.745 2794.230 145.575 ;
        RECT 5.330 137.305 2794.230 140.135 ;
        RECT 5.330 131.865 2794.230 134.695 ;
        RECT 5.330 126.425 2794.230 129.255 ;
        RECT 5.330 120.985 2794.230 123.815 ;
        RECT 5.330 115.545 2794.230 118.375 ;
        RECT 5.330 110.105 2794.230 112.935 ;
        RECT 5.330 104.665 2794.230 107.495 ;
        RECT 5.330 99.225 2794.230 102.055 ;
        RECT 5.330 93.785 2794.230 96.615 ;
        RECT 5.330 88.345 2794.230 91.175 ;
        RECT 5.330 82.905 2794.230 85.735 ;
        RECT 5.330 77.465 2794.230 80.295 ;
        RECT 5.330 72.025 2794.230 74.855 ;
        RECT 5.330 66.585 2794.230 69.415 ;
        RECT 5.330 61.145 2794.230 63.975 ;
        RECT 5.330 55.705 2794.230 58.535 ;
        RECT 5.330 50.265 2794.230 53.095 ;
        RECT 5.330 44.825 2794.230 47.655 ;
        RECT 5.330 39.385 2794.230 42.215 ;
        RECT 5.330 33.945 2794.230 36.775 ;
        RECT 5.330 28.505 2794.230 31.335 ;
        RECT 5.330 23.065 2794.230 25.895 ;
        RECT 5.330 17.625 2794.230 20.455 ;
        RECT 5.330 12.185 2794.230 15.015 ;
      LAYER li1 ;
        RECT 5.520 10.795 2794.040 1749.045 ;
      LAYER met1 ;
        RECT 5.520 0.720 2794.040 1749.200 ;
      LAYER met2 ;
        RECT 21.070 4.280 2787.410 1749.145 ;
        RECT 21.070 0.155 34.770 4.280 ;
        RECT 35.610 0.155 55.930 4.280 ;
        RECT 56.770 0.155 77.090 4.280 ;
        RECT 77.930 0.155 98.250 4.280 ;
        RECT 99.090 0.155 119.410 4.280 ;
        RECT 120.250 0.155 140.570 4.280 ;
        RECT 141.410 0.155 161.730 4.280 ;
        RECT 162.570 0.155 182.890 4.280 ;
        RECT 183.730 0.155 204.050 4.280 ;
        RECT 204.890 0.155 225.210 4.280 ;
        RECT 226.050 0.155 246.370 4.280 ;
        RECT 247.210 0.155 267.530 4.280 ;
        RECT 268.370 0.155 288.690 4.280 ;
        RECT 289.530 0.155 309.850 4.280 ;
        RECT 310.690 0.155 331.010 4.280 ;
        RECT 331.850 0.155 352.170 4.280 ;
        RECT 353.010 0.155 373.330 4.280 ;
        RECT 374.170 0.155 394.490 4.280 ;
        RECT 395.330 0.155 415.650 4.280 ;
        RECT 416.490 0.155 436.810 4.280 ;
        RECT 437.650 0.155 457.970 4.280 ;
        RECT 458.810 0.155 479.130 4.280 ;
        RECT 479.970 0.155 500.290 4.280 ;
        RECT 501.130 0.155 521.450 4.280 ;
        RECT 522.290 0.155 542.610 4.280 ;
        RECT 543.450 0.155 563.770 4.280 ;
        RECT 564.610 0.155 584.930 4.280 ;
        RECT 585.770 0.155 606.090 4.280 ;
        RECT 606.930 0.155 627.250 4.280 ;
        RECT 628.090 0.155 648.410 4.280 ;
        RECT 649.250 0.155 669.570 4.280 ;
        RECT 670.410 0.155 690.730 4.280 ;
        RECT 691.570 0.155 711.890 4.280 ;
        RECT 712.730 0.155 733.050 4.280 ;
        RECT 733.890 0.155 754.210 4.280 ;
        RECT 755.050 0.155 775.370 4.280 ;
        RECT 776.210 0.155 796.530 4.280 ;
        RECT 797.370 0.155 817.690 4.280 ;
        RECT 818.530 0.155 838.850 4.280 ;
        RECT 839.690 0.155 860.010 4.280 ;
        RECT 860.850 0.155 881.170 4.280 ;
        RECT 882.010 0.155 902.330 4.280 ;
        RECT 903.170 0.155 923.490 4.280 ;
        RECT 924.330 0.155 944.650 4.280 ;
        RECT 945.490 0.155 965.810 4.280 ;
        RECT 966.650 0.155 986.970 4.280 ;
        RECT 987.810 0.155 1008.130 4.280 ;
        RECT 1008.970 0.155 1029.290 4.280 ;
        RECT 1030.130 0.155 1050.450 4.280 ;
        RECT 1051.290 0.155 1071.610 4.280 ;
        RECT 1072.450 0.155 1092.770 4.280 ;
        RECT 1093.610 0.155 1113.930 4.280 ;
        RECT 1114.770 0.155 1135.090 4.280 ;
        RECT 1135.930 0.155 1156.250 4.280 ;
        RECT 1157.090 0.155 1177.410 4.280 ;
        RECT 1178.250 0.155 1198.570 4.280 ;
        RECT 1199.410 0.155 1219.730 4.280 ;
        RECT 1220.570 0.155 1240.890 4.280 ;
        RECT 1241.730 0.155 1262.050 4.280 ;
        RECT 1262.890 0.155 1283.210 4.280 ;
        RECT 1284.050 0.155 1304.370 4.280 ;
        RECT 1305.210 0.155 1325.530 4.280 ;
        RECT 1326.370 0.155 1346.690 4.280 ;
        RECT 1347.530 0.155 1367.850 4.280 ;
        RECT 1368.690 0.155 1389.010 4.280 ;
        RECT 1389.850 0.155 1410.170 4.280 ;
        RECT 1411.010 0.155 1431.330 4.280 ;
        RECT 1432.170 0.155 1452.490 4.280 ;
        RECT 1453.330 0.155 1473.650 4.280 ;
        RECT 1474.490 0.155 1494.810 4.280 ;
        RECT 1495.650 0.155 1515.970 4.280 ;
        RECT 1516.810 0.155 1537.130 4.280 ;
        RECT 1537.970 0.155 1558.290 4.280 ;
        RECT 1559.130 0.155 1579.450 4.280 ;
        RECT 1580.290 0.155 1600.610 4.280 ;
        RECT 1601.450 0.155 1621.770 4.280 ;
        RECT 1622.610 0.155 1642.930 4.280 ;
        RECT 1643.770 0.155 1664.090 4.280 ;
        RECT 1664.930 0.155 1685.250 4.280 ;
        RECT 1686.090 0.155 1706.410 4.280 ;
        RECT 1707.250 0.155 1727.570 4.280 ;
        RECT 1728.410 0.155 1748.730 4.280 ;
        RECT 1749.570 0.155 1769.890 4.280 ;
        RECT 1770.730 0.155 1791.050 4.280 ;
        RECT 1791.890 0.155 1812.210 4.280 ;
        RECT 1813.050 0.155 1833.370 4.280 ;
        RECT 1834.210 0.155 1854.530 4.280 ;
        RECT 1855.370 0.155 1875.690 4.280 ;
        RECT 1876.530 0.155 1896.850 4.280 ;
        RECT 1897.690 0.155 1918.010 4.280 ;
        RECT 1918.850 0.155 1939.170 4.280 ;
        RECT 1940.010 0.155 1960.330 4.280 ;
        RECT 1961.170 0.155 1981.490 4.280 ;
        RECT 1982.330 0.155 2002.650 4.280 ;
        RECT 2003.490 0.155 2023.810 4.280 ;
        RECT 2024.650 0.155 2044.970 4.280 ;
        RECT 2045.810 0.155 2066.130 4.280 ;
        RECT 2066.970 0.155 2087.290 4.280 ;
        RECT 2088.130 0.155 2108.450 4.280 ;
        RECT 2109.290 0.155 2129.610 4.280 ;
        RECT 2130.450 0.155 2150.770 4.280 ;
        RECT 2151.610 0.155 2171.930 4.280 ;
        RECT 2172.770 0.155 2193.090 4.280 ;
        RECT 2193.930 0.155 2214.250 4.280 ;
        RECT 2215.090 0.155 2235.410 4.280 ;
        RECT 2236.250 0.155 2256.570 4.280 ;
        RECT 2257.410 0.155 2277.730 4.280 ;
        RECT 2278.570 0.155 2298.890 4.280 ;
        RECT 2299.730 0.155 2320.050 4.280 ;
        RECT 2320.890 0.155 2341.210 4.280 ;
        RECT 2342.050 0.155 2362.370 4.280 ;
        RECT 2363.210 0.155 2383.530 4.280 ;
        RECT 2384.370 0.155 2404.690 4.280 ;
        RECT 2405.530 0.155 2425.850 4.280 ;
        RECT 2426.690 0.155 2447.010 4.280 ;
        RECT 2447.850 0.155 2468.170 4.280 ;
        RECT 2469.010 0.155 2489.330 4.280 ;
        RECT 2490.170 0.155 2510.490 4.280 ;
        RECT 2511.330 0.155 2531.650 4.280 ;
        RECT 2532.490 0.155 2552.810 4.280 ;
        RECT 2553.650 0.155 2573.970 4.280 ;
        RECT 2574.810 0.155 2595.130 4.280 ;
        RECT 2595.970 0.155 2616.290 4.280 ;
        RECT 2617.130 0.155 2637.450 4.280 ;
        RECT 2638.290 0.155 2658.610 4.280 ;
        RECT 2659.450 0.155 2679.770 4.280 ;
        RECT 2680.610 0.155 2700.930 4.280 ;
        RECT 2701.770 0.155 2722.090 4.280 ;
        RECT 2722.930 0.155 2743.250 4.280 ;
        RECT 2744.090 0.155 2764.410 4.280 ;
        RECT 2765.250 0.155 2787.410 4.280 ;
      LAYER met3 ;
        RECT 21.050 0.175 2787.430 1749.125 ;
      LAYER met4 ;
        RECT 958.015 10.240 1019.040 148.065 ;
        RECT 1021.440 10.240 1095.840 148.065 ;
        RECT 1098.240 10.240 1172.640 148.065 ;
        RECT 1175.040 10.240 1249.440 148.065 ;
        RECT 1251.840 10.240 1326.240 148.065 ;
        RECT 1328.640 10.240 1390.745 148.065 ;
        RECT 958.015 0.175 1390.745 10.240 ;
  END
END user_proj_example
END LIBRARY

