module __masc__execute (
	clk,
	instruction,
	rs1,
	rs2,
	bs,
	valid,
	out
);
	input wire clk;
	input wire [31:0] instruction;
	input wire [31:0] rs1;
	input wire [31:0] rs2;
	input wire [7:0] bs;
	input wire valid;
	output wire [32:0] out;
	wire [2047:0] inv_sbox__1;
	assign inv_sbox__1 = 2048'h52096ad53036a538bf40a39e81f3d7fb7ce339829b2fff87348e4344c4dee9cb547b9432a6c2233dee4c950b42fac34e082ea16628d924b2765ba2496d8bd12572f8f66486689816d4a45ccc5d65b6926c704850fdedb9da5e154657a78d9d8490d8ab008cbcd30af7e45805b8b34506d02c1e8fca3f0f02c1afbd0301138a6b3a9111414f67dcea97f2cfcef0b4e67396ac7422e7ad3585e2f937e81c75df6e47f11a711d29c5896fb7620eaa18be1bfc563e4bc6d279209adbc0fe78cd5af41fdda8338807c731b11210592780ec5f60517fa919b54a0d2de57a9f93c99cefa0e03b4dae2af5b0c8ebbb3c83539961172b047eba77d626e169146355210c7d;
	reg [31:0] p0_instruction;
	reg [31:0] p0_rs1;
	reg [31:0] p0_rs2;
	reg [7:0] p0_bs;
	reg p0_valid;
	always @(posedge clk) begin
		p0_instruction <= instruction;
		p0_rs1 <= rs1;
		p0_rs2 <= rs2;
		p0_bs <= bs;
		p0_valid <= valid;
	end
	wire [4:0] p1_bit_slice_13185_comb;
	wire [2:0] p1_literal_13186_comb;
	wire [1:0] p1_bit_slice_13190_comb;
	wire [2:0] p1_literal_13191_comb;
	wire [7:0] p1_shamt__2_comb;
	wire [4:0] p1_concat_13192_comb;
	wire [31:0] p1_literal_13243_comb;
	wire [31:0] p1_shrl_13188_comb;
	wire [31:0] p1_shrl_13193_comb;
	wire [31:0] p1_literal_13195_comb;
	wire [31:0] p1_literal_13196_comb;
	wire [31:0] p1_literal_13197_comb;
	wire [31:0] p1_literal_13198_comb;
	wire [31:0] p1_literal_13199_comb;
	wire [31:0] p1_literal_13200_comb;
	wire [31:0] p1_literal_13201_comb;
	wire [31:0] p1_literal_13202_comb;
	wire [31:0] p1_literal_13205_comb;
	wire [31:0] p1_literal_13206_comb;
	wire [31:0] p1_literal_13207_comb;
	wire [31:0] p1_literal_13208_comb;
	wire [31:0] p1_literal_13209_comb;
	wire [31:0] p1_literal_13210_comb;
	wire [31:0] p1_literal_13211_comb;
	wire [31:0] p1_literal_13212_comb;
	wire [31:0] p1_literal_13213_comb;
	wire [31:0] p1_literal_13216_comb;
	wire [31:0] p1_literal_13217_comb;
	wire [31:0] p1_literal_13218_comb;
	wire [31:0] p1_literal_13219_comb;
	wire [31:0] p1_literal_13220_comb;
	wire [31:0] p1_literal_13221_comb;
	wire [31:0] p1_literal_13222_comb;
	wire p1_ult_13244_comb;
	wire [7:0] p1_si__1_comb;
	wire [7:0] p1_si__2_comb;
	wire p1_eq_13203_comb;
	wire p1_eq_13204_comb;
	wire p1_eq_13214_comb;
	wire p1_eq_13215_comb;
	wire p1_eq_13223_comb;
	wire p1_eq_13224_comb;
	wire p1_eq_13225_comb;
	wire p1_eq_13226_comb;
	wire p1_eq_13227_comb;
	wire p1_eq_13228_comb;
	wire p1_eq_13229_comb;
	wire p1_eq_13230_comb;
	wire p1_eq_13231_comb;
	wire p1_eq_13232_comb;
	wire p1_eq_13233_comb;
	wire p1_eq_13234_comb;
	wire p1_eq_13235_comb;
	wire p1_eq_13236_comb;
	wire p1_eq_13237_comb;
	wire p1_eq_13238_comb;
	wire p1_eq_13239_comb;
	wire p1_eq_13240_comb;
	wire p1_eq_13241_comb;
	wire p1_eq_13242_comb;
	wire p1_and_13245_comb;
	assign p1_bit_slice_13185_comb = p0_bs[4:0];
	assign p1_literal_13186_comb = 3'h0;
	assign p1_bit_slice_13190_comb = p0_bs[1:0];
	assign p1_literal_13191_comb = 3'h0;
	assign p1_shamt__2_comb = {p1_bit_slice_13185_comb, p1_literal_13186_comb};
	assign p1_concat_13192_comb = {p1_bit_slice_13190_comb, p1_literal_13191_comb};
	assign p1_literal_13243_comb = 32'h00000018;
	assign p1_shrl_13188_comb = (p1_shamt__2_comb >= 8'h20 ? 32'h00000000 : p0_rs2 >> p1_shamt__2_comb);
	assign p1_shrl_13193_comb = p0_rs2 >> p1_concat_13192_comb;
	assign p1_literal_13195_comb = 32'h00000006;
	assign p1_literal_13196_comb = 32'h00000007;
	assign p1_literal_13197_comb = 32'h0000000a;
	assign p1_literal_13198_comb = 32'h0000000b;
	assign p1_literal_13199_comb = 32'h00000011;
	assign p1_literal_13200_comb = 32'h00000013;
	assign p1_literal_13201_comb = 32'h00000009;
	assign p1_literal_13202_comb = 32'h00000014;
	assign p1_literal_13205_comb = 32'h00000017;
	assign p1_literal_13206_comb = 32'h00000016;
	assign p1_literal_13207_comb = 32'h00000015;
	assign p1_literal_13208_comb = 32'h00000012;
	assign p1_literal_13209_comb = 32'h00000010;
	assign p1_literal_13210_comb = 32'h0000000f;
	assign p1_literal_13211_comb = 32'h0000000e;
	assign p1_literal_13212_comb = 32'h0000000d;
	assign p1_literal_13213_comb = 32'h0000000c;
	assign p1_literal_13216_comb = 32'h00000008;
	assign p1_literal_13217_comb = 32'h00000005;
	assign p1_literal_13218_comb = 32'h00000004;
	assign p1_literal_13219_comb = 32'h00000003;
	assign p1_literal_13220_comb = 32'h00000002;
	assign p1_literal_13221_comb = 32'h00000001;
	assign p1_literal_13222_comb = 32'h00000000;
	assign p1_ult_13244_comb = p0_instruction < p1_literal_13243_comb;
	assign p1_si__1_comb = p1_shrl_13188_comb[7:0];
	assign p1_si__2_comb = p1_shrl_13193_comb[7:0];
	assign p1_eq_13203_comb = p0_instruction == p1_literal_13195_comb;
	assign p1_eq_13204_comb = p0_instruction == p1_literal_13196_comb;
	assign p1_eq_13214_comb = p0_instruction == p1_literal_13197_comb;
	assign p1_eq_13215_comb = p0_instruction == p1_literal_13198_comb;
	assign p1_eq_13223_comb = p0_instruction == p1_literal_13199_comb;
	assign p1_eq_13224_comb = p0_instruction == p1_literal_13200_comb;
	assign p1_eq_13225_comb = p0_instruction == p1_literal_13201_comb;
	assign p1_eq_13226_comb = p0_instruction == p1_literal_13202_comb;
	assign p1_eq_13227_comb = p0_instruction == p1_literal_13205_comb;
	assign p1_eq_13228_comb = p0_instruction == p1_literal_13206_comb;
	assign p1_eq_13229_comb = p0_instruction == p1_literal_13207_comb;
	assign p1_eq_13230_comb = p0_instruction == p1_literal_13208_comb;
	assign p1_eq_13231_comb = p0_instruction == p1_literal_13209_comb;
	assign p1_eq_13232_comb = p0_instruction == p1_literal_13210_comb;
	assign p1_eq_13233_comb = p0_instruction == p1_literal_13211_comb;
	assign p1_eq_13234_comb = p0_instruction == p1_literal_13212_comb;
	assign p1_eq_13235_comb = p0_instruction == p1_literal_13213_comb;
	assign p1_eq_13236_comb = p0_instruction == p1_literal_13216_comb;
	assign p1_eq_13237_comb = p0_instruction == p1_literal_13217_comb;
	assign p1_eq_13238_comb = p0_instruction == p1_literal_13218_comb;
	assign p1_eq_13239_comb = p0_instruction == p1_literal_13219_comb;
	assign p1_eq_13240_comb = p0_instruction == p1_literal_13220_comb;
	assign p1_eq_13241_comb = p0_instruction == p1_literal_13221_comb;
	assign p1_eq_13242_comb = p0_instruction == p1_literal_13222_comb;
	assign p1_and_13245_comb = p0_valid & p1_ult_13244_comb;
	reg [31:0] p1_rs1;
	reg [31:0] p1_rs2;
	reg p1_valid;
	reg [7:0] p1_si__1;
	reg [1:0] p1_bit_slice_13190;
	reg [4:0] p1_concat_13192;
	reg [7:0] p1_si__2;
	reg p1_eq_13203;
	reg p1_eq_13204;
	reg p1_eq_13214;
	reg p1_eq_13215;
	reg p1_eq_13223;
	reg p1_eq_13224;
	reg p1_eq_13225;
	reg p1_eq_13226;
	reg p1_eq_13227;
	reg p1_eq_13228;
	reg p1_eq_13229;
	reg p1_eq_13230;
	reg p1_eq_13231;
	reg p1_eq_13232;
	reg p1_eq_13233;
	reg p1_eq_13234;
	reg p1_eq_13235;
	reg p1_eq_13236;
	reg p1_eq_13237;
	reg p1_eq_13238;
	reg p1_eq_13239;
	reg p1_eq_13240;
	reg p1_eq_13241;
	reg p1_eq_13242;
	reg p1_and_13245;
	always @(posedge clk) begin
		p1_rs1 <= p0_rs1;
		p1_rs2 <= p0_rs2;
		p1_valid <= p0_valid;
		p1_si__1 <= p1_si__1_comb;
		p1_bit_slice_13190 <= p1_bit_slice_13190_comb;
		p1_concat_13192 <= p1_concat_13192_comb;
		p1_si__2 <= p1_si__2_comb;
		p1_eq_13203 <= p1_eq_13203_comb;
		p1_eq_13204 <= p1_eq_13204_comb;
		p1_eq_13214 <= p1_eq_13214_comb;
		p1_eq_13215 <= p1_eq_13215_comb;
		p1_eq_13223 <= p1_eq_13223_comb;
		p1_eq_13224 <= p1_eq_13224_comb;
		p1_eq_13225 <= p1_eq_13225_comb;
		p1_eq_13226 <= p1_eq_13226_comb;
		p1_eq_13227 <= p1_eq_13227_comb;
		p1_eq_13228 <= p1_eq_13228_comb;
		p1_eq_13229 <= p1_eq_13229_comb;
		p1_eq_13230 <= p1_eq_13230_comb;
		p1_eq_13231 <= p1_eq_13231_comb;
		p1_eq_13232 <= p1_eq_13232_comb;
		p1_eq_13233 <= p1_eq_13233_comb;
		p1_eq_13234 <= p1_eq_13234_comb;
		p1_eq_13235 <= p1_eq_13235_comb;
		p1_eq_13236 <= p1_eq_13236_comb;
		p1_eq_13237 <= p1_eq_13237_comb;
		p1_eq_13238 <= p1_eq_13238_comb;
		p1_eq_13239 <= p1_eq_13239_comb;
		p1_eq_13240 <= p1_eq_13240_comb;
		p1_eq_13241 <= p1_eq_13241_comb;
		p1_eq_13242 <= p1_eq_13242_comb;
		p1_and_13245 <= p1_and_13245_comb;
	end
	wire [7:0] p2_so__1_comb;
	wire [7:0] p2_sbox_inv_val_comb;
	assign p2_so__1_comb = inv_sbox__1[(255 - p1_si__1) * 8+:8];
	assign p2_sbox_inv_val_comb = inv_sbox__1[(255 - p1_si__2) * 8+:8];
	reg [31:0] p2_rs1;
	reg [31:0] p2_rs2;
	reg p2_valid;
	reg [7:0] p2_so__1;
	reg [1:0] p2_bit_slice_13190;
	reg [4:0] p2_concat_13192;
	reg [7:0] p2_sbox_inv_val;
	reg p2_eq_13203;
	reg p2_eq_13204;
	reg p2_eq_13214;
	reg p2_eq_13215;
	reg p2_eq_13223;
	reg p2_eq_13224;
	reg p2_eq_13225;
	reg p2_eq_13226;
	reg p2_eq_13227;
	reg p2_eq_13228;
	reg p2_eq_13229;
	reg p2_eq_13230;
	reg p2_eq_13231;
	reg p2_eq_13232;
	reg p2_eq_13233;
	reg p2_eq_13234;
	reg p2_eq_13235;
	reg p2_eq_13236;
	reg p2_eq_13237;
	reg p2_eq_13238;
	reg p2_eq_13239;
	reg p2_eq_13240;
	reg p2_eq_13241;
	reg p2_eq_13242;
	reg p2_and_13245;
	always @(posedge clk) begin
		p2_rs1 <= p1_rs1;
		p2_rs2 <= p1_rs2;
		p2_valid <= p1_valid;
		p2_so__1 <= p2_so__1_comb;
		p2_bit_slice_13190 <= p1_bit_slice_13190;
		p2_concat_13192 <= p1_concat_13192;
		p2_sbox_inv_val <= p2_sbox_inv_val_comb;
		p2_eq_13203 <= p1_eq_13203;
		p2_eq_13204 <= p1_eq_13204;
		p2_eq_13214 <= p1_eq_13214;
		p2_eq_13215 <= p1_eq_13215;
		p2_eq_13223 <= p1_eq_13223;
		p2_eq_13224 <= p1_eq_13224;
		p2_eq_13225 <= p1_eq_13225;
		p2_eq_13226 <= p1_eq_13226;
		p2_eq_13227 <= p1_eq_13227;
		p2_eq_13228 <= p1_eq_13228;
		p2_eq_13229 <= p1_eq_13229;
		p2_eq_13230 <= p1_eq_13230;
		p2_eq_13231 <= p1_eq_13231;
		p2_eq_13232 <= p1_eq_13232;
		p2_eq_13233 <= p1_eq_13233;
		p2_eq_13234 <= p1_eq_13234;
		p2_eq_13235 <= p1_eq_13235;
		p2_eq_13236 <= p1_eq_13236;
		p2_eq_13237 <= p1_eq_13237;
		p2_eq_13238 <= p1_eq_13238;
		p2_eq_13239 <= p1_eq_13239;
		p2_eq_13240 <= p1_eq_13240;
		p2_eq_13241 <= p1_eq_13241;
		p2_eq_13242 <= p1_eq_13242;
		p2_and_13245 <= p1_and_13245;
	end
	wire p3_bit_slice_13377_comb;
	wire [6:0] p3_bit_slice_13378_comb;
	wire p3_literal_13379_comb;
	wire [7:0] p3_sign_ext_13380_comb;
	wire [7:0] p3_literal_13381_comb;
	wire [7:0] p3_xshifted_comb;
	wire [7:0] p3_conditional_xor__1_comb;
	wire [7:0] p3_term_2_comb;
	wire p3_bit_slice_13385_comb;
	wire [6:0] p3_bit_slice_13386_comb;
	wire p3_literal_13387_comb;
	wire [7:0] p3_sign_ext_13388_comb;
	wire [7:0] p3_literal_13389_comb;
	wire [7:0] p3_xshifted__1_comb;
	wire [7:0] p3_conditional_xor__2_comb;
	wire [7:0] p3_term_3__1_comb;
	wire p3_bit_slice_13393_comb;
	wire [6:0] p3_bit_slice_13394_comb;
	wire p3_literal_13395_comb;
	wire [7:0] p3_sign_ext_13396_comb;
	wire [7:0] p3_literal_13397_comb;
	wire [7:0] p3_xshifted__2_comb;
	wire [7:0] p3_conditional_xor__3_comb;
	wire p3_literal_13400_comb;
	wire [2:0] p3_literal_13401_comb;
	wire [7:0] p3_term_4_comb;
	wire p3_literal_13403_comb;
	wire [4:0] p3_bit_slice_13404_comb;
	wire [5:0] p3_literal_13405_comb;
	wire [5:0] p3_concat_13406_comb;
	wire [7:0] p3_xor_13407_comb;
	wire [7:0] p3_xor_13408_comb;
	wire [7:0] p3_xor_13409_comb;
	wire [7:0] p3_xor_13410_comb;
	wire [5:0] p3_literal_13411_comb;
	wire [5:0] p3_concat_13412_comb;
	wire [31:0] p3_literal_13413_comb;
	wire [5:0] p3_sub_13414_comb;
	wire [31:0] p3_mixed_comb;
	wire [5:0] p3_sub_13416_comb;
	wire [31:0] p3_sub_13417_comb;
	assign p3_bit_slice_13377_comb = p2_so__1[7];
	assign p3_bit_slice_13378_comb = p2_so__1[6:0];
	assign p3_literal_13379_comb = 1'h0;
	assign p3_sign_ext_13380_comb = {8 {p3_bit_slice_13377_comb}};
	assign p3_literal_13381_comb = 8'h1b;
	assign p3_xshifted_comb = {p3_bit_slice_13378_comb, p3_literal_13379_comb};
	assign p3_conditional_xor__1_comb = p3_sign_ext_13380_comb & p3_literal_13381_comb;
	assign p3_term_2_comb = p3_xshifted_comb ^ p3_conditional_xor__1_comb;
	assign p3_bit_slice_13385_comb = p3_term_2_comb[7];
	assign p3_bit_slice_13386_comb = p3_term_2_comb[6:0];
	assign p3_literal_13387_comb = 1'h0;
	assign p3_sign_ext_13388_comb = {8 {p3_bit_slice_13385_comb}};
	assign p3_literal_13389_comb = 8'h1b;
	assign p3_xshifted__1_comb = {p3_bit_slice_13386_comb, p3_literal_13387_comb};
	assign p3_conditional_xor__2_comb = p3_sign_ext_13388_comb & p3_literal_13389_comb;
	assign p3_term_3__1_comb = p3_xshifted__1_comb ^ p3_conditional_xor__2_comb;
	assign p3_bit_slice_13393_comb = p3_term_3__1_comb[7];
	assign p3_bit_slice_13394_comb = p3_term_3__1_comb[6:0];
	assign p3_literal_13395_comb = 1'h0;
	assign p3_sign_ext_13396_comb = {8 {p3_bit_slice_13393_comb}};
	assign p3_literal_13397_comb = 8'h1b;
	assign p3_xshifted__2_comb = {p3_bit_slice_13394_comb, p3_literal_13395_comb};
	assign p3_conditional_xor__3_comb = p3_sign_ext_13396_comb & p3_literal_13397_comb;
	assign p3_literal_13400_comb = 1'h0;
	assign p3_literal_13401_comb = 3'h0;
	assign p3_term_4_comb = p3_xshifted__2_comb ^ p3_conditional_xor__3_comb;
	assign p3_literal_13403_comb = 1'h0;
	assign p3_bit_slice_13404_comb = p2_rs2[4:0];
	assign p3_literal_13405_comb = 6'h20;
	assign p3_concat_13406_comb = {p3_literal_13400_comb, p2_bit_slice_13190, p3_literal_13401_comb};
	assign p3_xor_13407_comb = (p2_so__1 ^ p3_term_2_comb) ^ p3_term_4_comb;
	assign p3_xor_13408_comb = (p2_so__1 ^ p3_term_3__1_comb) ^ p3_term_4_comb;
	assign p3_xor_13409_comb = p2_so__1 ^ p3_term_4_comb;
	assign p3_xor_13410_comb = (p3_term_2_comb ^ p3_term_3__1_comb) ^ p3_term_4_comb;
	assign p3_literal_13411_comb = 6'h20;
	assign p3_concat_13412_comb = {p3_literal_13403_comb, p3_bit_slice_13404_comb};
	assign p3_literal_13413_comb = 32'h00000020;
	assign p3_sub_13414_comb = p3_literal_13405_comb - p3_concat_13406_comb;
	assign p3_mixed_comb = {p3_xor_13407_comb, p3_xor_13408_comb, p3_xor_13409_comb, p3_xor_13410_comb};
	assign p3_sub_13416_comb = p3_literal_13411_comb - p3_concat_13412_comb;
	assign p3_sub_13417_comb = p3_literal_13413_comb - p2_rs2;
	reg [31:0] p3_rs1;
	reg [31:0] p3_rs2;
	reg p3_valid;
	reg [4:0] p3_concat_13192;
	reg [4:0] p3_bit_slice_13404;
	reg [7:0] p3_sbox_inv_val;
	reg [5:0] p3_sub_13414;
	reg [31:0] p3_mixed;
	reg [5:0] p3_sub_13416;
	reg [31:0] p3_sub_13417;
	reg p3_eq_13203;
	reg p3_eq_13204;
	reg p3_eq_13214;
	reg p3_eq_13215;
	reg p3_eq_13223;
	reg p3_eq_13224;
	reg p3_eq_13225;
	reg p3_eq_13226;
	reg p3_eq_13227;
	reg p3_eq_13228;
	reg p3_eq_13229;
	reg p3_eq_13230;
	reg p3_eq_13231;
	reg p3_eq_13232;
	reg p3_eq_13233;
	reg p3_eq_13234;
	reg p3_eq_13235;
	reg p3_eq_13236;
	reg p3_eq_13237;
	reg p3_eq_13238;
	reg p3_eq_13239;
	reg p3_eq_13240;
	reg p3_eq_13241;
	reg p3_eq_13242;
	reg p3_and_13245;
	always @(posedge clk) begin
		p3_rs1 <= p2_rs1;
		p3_rs2 <= p2_rs2;
		p3_valid <= p2_valid;
		p3_concat_13192 <= p2_concat_13192;
		p3_bit_slice_13404 <= p3_bit_slice_13404_comb;
		p3_sbox_inv_val <= p2_sbox_inv_val;
		p3_sub_13414 <= p3_sub_13414_comb;
		p3_mixed <= p3_mixed_comb;
		p3_sub_13416 <= p3_sub_13416_comb;
		p3_sub_13417 <= p3_sub_13417_comb;
		p3_eq_13203 <= p2_eq_13203;
		p3_eq_13204 <= p2_eq_13204;
		p3_eq_13214 <= p2_eq_13214;
		p3_eq_13215 <= p2_eq_13215;
		p3_eq_13223 <= p2_eq_13223;
		p3_eq_13224 <= p2_eq_13224;
		p3_eq_13225 <= p2_eq_13225;
		p3_eq_13226 <= p2_eq_13226;
		p3_eq_13227 <= p2_eq_13227;
		p3_eq_13228 <= p2_eq_13228;
		p3_eq_13229 <= p2_eq_13229;
		p3_eq_13230 <= p2_eq_13230;
		p3_eq_13231 <= p2_eq_13231;
		p3_eq_13232 <= p2_eq_13232;
		p3_eq_13233 <= p2_eq_13233;
		p3_eq_13234 <= p2_eq_13234;
		p3_eq_13235 <= p2_eq_13235;
		p3_eq_13236 <= p2_eq_13236;
		p3_eq_13237 <= p2_eq_13237;
		p3_eq_13238 <= p2_eq_13238;
		p3_eq_13239 <= p2_eq_13239;
		p3_eq_13240 <= p2_eq_13240;
		p3_eq_13241 <= p2_eq_13241;
		p3_eq_13242 <= p2_eq_13242;
		p3_and_13245 <= p2_and_13245;
	end
	wire [23:0] p4_literal_13488_comb;
	wire [31:0] p4_so__2_comb;
	wire [31:0] p4_shll_13490_comb;
	wire [31:0] p4_shrl_13491_comb;
	wire [31:0] p4_shll_13492_comb;
	wire [31:0] p4_shrl_13493_comb;
	wire [31:0] p4_shrl_13494_comb;
	wire [31:0] p4_shll_13495_comb;
	wire [31:0] p4_shll_13496_comb;
	wire [31:0] p4_shrl_13497_comb;
	wire [31:0] p4_shrl_13498_comb;
	wire [31:0] p4_shll_13499_comb;
	assign p4_literal_13488_comb = 24'h000000;
	assign p4_so__2_comb = {p4_literal_13488_comb, p3_sbox_inv_val};
	assign p4_shll_13490_comb = p4_so__2_comb << p3_concat_13192;
	assign p4_shrl_13491_comb = (p3_sub_13414 >= 6'h20 ? 32'h00000000 : p4_so__2_comb >> p3_sub_13414);
	assign p4_shll_13492_comb = p3_mixed << p3_concat_13192;
	assign p4_shrl_13493_comb = (p3_sub_13414 >= 6'h20 ? 32'h00000000 : p3_mixed >> p3_sub_13414);
	assign p4_shrl_13494_comb = p3_rs1 >> p3_bit_slice_13404;
	assign p4_shll_13495_comb = (p3_sub_13416 >= 6'h20 ? 32'h00000000 : p3_rs1 << p3_sub_13416);
	assign p4_shll_13496_comb = p3_rs1 << p3_bit_slice_13404;
	assign p4_shrl_13497_comb = (p3_sub_13416 >= 6'h20 ? 32'h00000000 : p3_rs1 >> p3_sub_13416);
	assign p4_shrl_13498_comb = (p3_rs2 >= 32'h00000020 ? 32'h00000000 : p3_rs1 >> p3_rs2);
	assign p4_shll_13499_comb = (p3_sub_13417 >= 32'h00000020 ? 32'h00000000 : p3_rs1 << p3_sub_13417);
	reg [31:0] p4_rs1;
	reg [31:0] p4_rs2;
	reg p4_valid;
	reg [31:0] p4_shll_13490;
	reg [31:0] p4_shrl_13491;
	reg [31:0] p4_shll_13492;
	reg [31:0] p4_shrl_13493;
	reg p4_eq_13203;
	reg p4_eq_13204;
	reg p4_eq_13214;
	reg p4_eq_13215;
	reg [31:0] p4_shrl_13494;
	reg [31:0] p4_shll_13495;
	reg [31:0] p4_shll_13496;
	reg [31:0] p4_shrl_13497;
	reg [31:0] p4_shrl_13498;
	reg [31:0] p4_shll_13499;
	reg p4_eq_13223;
	reg p4_eq_13224;
	reg p4_eq_13225;
	reg p4_eq_13226;
	reg p4_eq_13227;
	reg p4_eq_13228;
	reg p4_eq_13229;
	reg p4_eq_13230;
	reg p4_eq_13231;
	reg p4_eq_13232;
	reg p4_eq_13233;
	reg p4_eq_13234;
	reg p4_eq_13235;
	reg p4_eq_13236;
	reg p4_eq_13237;
	reg p4_eq_13238;
	reg p4_eq_13239;
	reg p4_eq_13240;
	reg p4_eq_13241;
	reg p4_eq_13242;
	reg p4_and_13245;
	always @(posedge clk) begin
		p4_rs1 <= p3_rs1;
		p4_rs2 <= p3_rs2;
		p4_valid <= p3_valid;
		p4_shll_13490 <= p4_shll_13490_comb;
		p4_shrl_13491 <= p4_shrl_13491_comb;
		p4_shll_13492 <= p4_shll_13492_comb;
		p4_shrl_13493 <= p4_shrl_13493_comb;
		p4_eq_13203 <= p3_eq_13203;
		p4_eq_13204 <= p3_eq_13204;
		p4_eq_13214 <= p3_eq_13214;
		p4_eq_13215 <= p3_eq_13215;
		p4_shrl_13494 <= p4_shrl_13494_comb;
		p4_shll_13495 <= p4_shll_13495_comb;
		p4_shll_13496 <= p4_shll_13496_comb;
		p4_shrl_13497 <= p4_shrl_13497_comb;
		p4_shrl_13498 <= p4_shrl_13498_comb;
		p4_shll_13499 <= p4_shll_13499_comb;
		p4_eq_13223 <= p3_eq_13223;
		p4_eq_13224 <= p3_eq_13224;
		p4_eq_13225 <= p3_eq_13225;
		p4_eq_13226 <= p3_eq_13226;
		p4_eq_13227 <= p3_eq_13227;
		p4_eq_13228 <= p3_eq_13228;
		p4_eq_13229 <= p3_eq_13229;
		p4_eq_13230 <= p3_eq_13230;
		p4_eq_13231 <= p3_eq_13231;
		p4_eq_13232 <= p3_eq_13232;
		p4_eq_13233 <= p3_eq_13233;
		p4_eq_13234 <= p3_eq_13234;
		p4_eq_13235 <= p3_eq_13235;
		p4_eq_13236 <= p3_eq_13236;
		p4_eq_13237 <= p3_eq_13237;
		p4_eq_13238 <= p3_eq_13238;
		p4_eq_13239 <= p3_eq_13239;
		p4_eq_13240 <= p3_eq_13240;
		p4_eq_13241 <= p3_eq_13241;
		p4_eq_13242 <= p3_eq_13242;
		p4_and_13245 <= p3_and_13245;
	end
	wire p5_rotation_1__6_comb;
	wire [30:0] p5_rotation_1__5_comb;
	wire [7:0] p5_byte0__1_comb;
	wire [23:0] p5_rotation_2__5_comb;
	wire [27:0] p5_rotation_1__10_comb;
	wire [3:0] p5_rotation_1__9_comb;
	wire [1:0] p5_rotation_2__10_comb;
	wire [29:0] p5_rotation_2__9_comb;
	wire [6:0] p5_literal_13584_comb;
	wire [24:0] p5_rotation_3__3_comb;
	wire [31:0] p5_rotation_1__1_comb;
	wire [31:0] p5_rotation_2__1_comb;
	wire [31:0] p5_rotation_1__2_comb;
	wire [31:0] p5_rotation_2__2_comb;
	wire [6:0] p5_rotation_3__4_comb;
	wire [1:0] p5_bit_slice_13591_comb;
	wire [1:0] p5_bit_slice_13592_comb;
	wire [4:0] p5_bit_slice_13593_comb;
	wire [4:0] p5_bit_slice_13594_comb;
	wire [4:0] p5_bit_slice_13595_comb;
	wire [1:0] p5_bit_slice_13596_comb;
	wire [1:0] p5_bit_slice_13597_comb;
	wire [10:0] p5_bit_slice_13598_comb;
	wire [10:0] p5_bit_slice_13599_comb;
	wire [10:0] p5_bit_slice_13600_comb;
	wire [2:0] p5_bit_slice_13601_comb;
	wire [2:0] p5_bit_slice_13602_comb;
	wire [3:0] p5_bit_slice_13603_comb;
	wire [3:0] p5_bit_slice_13604_comb;
	wire [20:0] p5_bit_slice_13605_comb;
	wire [20:0] p5_bit_slice_13606_comb;
	wire [20:0] p5_bit_slice_13607_comb;
	wire [10:0] p5_bit_slice_13608_comb;
	wire [8:0] p5_bit_slice_13609_comb;
	wire [8:0] p5_bit_slice_13610_comb;
	wire [8:0] p5_bit_slice_13611_comb;
	wire [4:0] p5_bit_slice_13612_comb;
	wire [13:0] p5_bit_slice_13613_comb;
	wire [13:0] p5_rotate_18__1_comb;
	wire [13:0] p5_bit_slice_13615_comb;
	wire [9:0] p5_bit_slice_13616_comb;
	wire [9:0] p5_bit_slice_13617_comb;
	wire [6:0] p5_bit_slice_13618_comb;
	wire [6:0] p5_rotation_3__5_comb;
	wire [13:0] p5_bit_slice_13620_comb;
	wire [13:0] p5_bit_slice_13621_comb;
	wire [9:0] p5_bit_slice_13622_comb;
	wire [9:0] p5_bit_slice_13623_comb;
	wire [9:0] p5_rot_c__1_comb;
	wire [3:0] p5_bit_slice_13625_comb;
	wire [3:0] p5_bit_slice_13626_comb;
	wire [6:0] p5_bit_slice_13627_comb;
	wire [6:0] p5_bit_slice_13628_comb;
	wire [31:0] p5_not_13629_comb;
	wire [31:0] p5_xor_13630_comb;
	wire [31:0] p5_shift_1_comb;
	wire [31:0] p5_combined_1_comb;
	wire [31:0] p5_combined_2_comb;
	wire [5:0] p5_rotation_1__12_comb;
	wire [5:0] p5_bit_slice_13635_comb;
	wire [5:0] p5_bit_slice_13636_comb;
	wire [5:0] p5_bit_slice_13637_comb;
	wire [5:0] p5_bit_slice_13638_comb;
	wire [31:0] p5_combined_1__1_comb;
	wire [31:0] p5_combined_2__1_comb;
	wire [31:0] p5_rotation_3__1_comb;
	wire [5:0] p5_bit_slice_13642_comb;
	wire [5:0] p5_bit_slice_13643_comb;
	wire [31:0] p5_or_13644_comb;
	wire [31:0] p5_or_13645_comb;
	wire [1:0] p5_result__44_comb;
	wire [4:0] p5_result__43_comb;
	wire [1:0] p5_xor_13648_comb;
	wire [10:0] p5_xor_13649_comb;
	wire [2:0] p5_xor_13650_comb;
	wire [3:0] p5_xor_13651_comb;
	wire [20:0] p5_result__42_comb;
	wire [10:0] p5_xor_13653_comb;
	wire [12:0] p5_bit_slice_13654_comb;
	wire [12:0] p5_rotation_1__13_comb;
	wire [12:0] p5_bit_slice_13656_comb;
	wire [12:0] p5_bit_slice_13657_comb;
	wire [8:0] p5_xor_13658_comb;
	wire [4:0] p5_xor_13659_comb;
	wire [13:0] p5_xor_13660_comb;
	wire [9:0] p5_xor_13661_comb;
	wire [6:0] p5_xor_13662_comb;
	wire [13:0] p5_xor_13663_comb;
	wire [9:0] p5_xor_13664_comb;
	wire [9:0] p5_bit_slice_13665_comb;
	wire [12:0] p5_bit_slice_13666_comb;
	wire [3:0] p5_result__41_comb;
	wire [6:0] p5_xor_13668_comb;
	wire [2:0] p5_bit_slice_13669_comb;
	wire [2:0] p5_bit_slice_13670_comb;
	wire [2:0] p5_bit_slice_13671_comb;
	wire [2:0] p5_rotation_2__13_comb;
	wire p5_or_13673_comb;
	wire p5_or_13674_comb;
	wire [31:0] p5_or_13675_comb;
	wire [31:0] p5_or_13676_comb;
	wire [31:0] p5_or_13677_comb;
	wire [31:0] p5_nor_13678_comb;
	wire [31:0] p5_nand_13679_comb;
	wire [31:0] p5_not_13680_comb;
	wire [31:0] p5_xor_13681_comb;
	wire [5:0] p5_xor_13682_comb;
	wire [5:0] p5_xor_13683_comb;
	wire [31:0] p5_xor_13684_comb;
	wire [5:0] p5_result__4_comb;
	wire [5:0] p5_xor_13686_comb;
	wire [31:0] p5_result__7_comb;
	wire [31:0] p5_result__8_comb;
	wire p5_result__28_comb;
	wire p5_result__30_comb;
	wire p5_result__32_comb;
	wire p5_result__34_comb;
	wire p5_result__36_comb;
	wire p5_result__39_comb;
	wire p5_result__38_comb;
	wire p5_result__37_comb;
	wire p5_result__35_comb;
	wire p5_result__24_comb;
	wire p5_result__20_comb;
	wire p5_bit_slice_13700_comb;
	wire [3:0] p5_bit_slice_13701_comb;
	wire p5_bit_slice_13702_comb;
	wire [3:0] p5_bit_slice_13703_comb;
	wire [1:0] p5_bit_slice_13704_comb;
	wire [2:0] p5_bit_slice_13705_comb;
	wire p5_or_13706_comb;
	wire p5_result__40_comb;
	wire p5_result__33_comb;
	wire p5_result__16_comb;
	wire p5_result__12_comb;
	wire p5_bit_slice_13711_comb;
	wire p5_bit_slice_13712_comb;
	wire p5_bit_slice_13713_comb;
	wire p5_bit_slice_13714_comb;
	wire [12:0] p5_result__3_comb;
	wire [12:0] p5_xor_13716_comb;
	wire p5_or_13717_comb;
	wire p5_result__14_comb;
	wire p5_result__18_comb;
	wire p5_result__22_comb;
	wire p5_result__31_comb;
	wire p5_result__29_comb;
	wire p5_result__27_comb;
	wire p5_result__26_comb;
	wire p5_result__23_comb;
	wire p5_result__19_comb;
	wire p5_result__15_comb;
	wire [3:0] p5_bit_slice_13728_comb;
	wire [1:0] p5_bit_slice_13729_comb;
	wire [1:0] p5_bit_slice_13730_comb;
	wire [3:0] p5_bit_slice_13731_comb;
	wire p5_bit_slice_13732_comb;
	wire [4:0] p5_bit_slice_13733_comb;
	wire p5_or_13734_comb;
	wire p5_bit_slice_13735_comb;
	wire p5_literal_13736_comb;
	wire p5_bit_slice_13737_comb;
	wire p5_result__25_comb;
	wire p5_result__11_comb;
	wire p5_bit_slice_13740_comb;
	wire p5_bit_slice_13741_comb;
	wire [1:0] p5_bit_slice_13742_comb;
	wire [1:0] p5_bit_slice_13743_comb;
	wire p5_or_13744_comb;
	wire p5_result__21_comb;
	wire [2:0] p5_bit_slice_13746_comb;
	wire p5_bit_slice_13747_comb;
	wire [9:0] p5_result__2_comb;
	wire [12:0] p5_xor_13749_comb;
	wire p5_result__13_comb;
	wire p5_result__17_comb;
	wire [3:0] p5_bit_slice_13752_comb;
	wire p5_bit_slice_13753_comb;
	wire p5_bit_slice_13754_comb;
	wire [3:0] p5_bit_slice_13755_comb;
	wire p5_result__10_comb;
	wire [2:0] p5_result__5_comb;
	wire [2:0] p5_xor_13758_comb;
	wire p5_or_13759_comb;
	wire [21:0] p5_concat_13760_comb;
	wire p5_bit_slice_13761_comb;
	wire p5_bit_slice_13762_comb;
	wire p5_bit_slice_13763_comb;
	wire p5_bit_slice_13764_comb;
	wire p5_bit_slice_13765_comb;
	wire p5_bit_slice_13766_comb;
	wire p5_bit_slice_13767_comb;
	wire p5_bit_slice_13768_comb;
	wire p5_bit_slice_13769_comb;
	wire p5_bit_slice_13770_comb;
	wire p5_bit_slice_13771_comb;
	wire p5_bit_slice_13772_comb;
	wire p5_bit_slice_13773_comb;
	wire p5_bit_slice_13774_comb;
	wire p5_bit_slice_13775_comb;
	wire p5_bit_slice_13776_comb;
	wire p5_bit_slice_13777_comb;
	wire p5_bit_slice_13778_comb;
	wire p5_bit_slice_13779_comb;
	wire [22:0] p5_concat_13780_comb;
	wire [4:0] p5_bit_slice_13781_comb;
	wire [4:0] p5_bit_slice_13782_comb;
	wire [4:0] p5_bit_slice_13783_comb;
	wire [4:0] p5_bit_slice_13784_comb;
	wire [4:0] p5_bit_slice_13785_comb;
	wire [4:0] p5_bit_slice_13786_comb;
	wire [4:0] p5_bit_slice_13787_comb;
	wire [4:0] p5_concat_13788_comb;
	wire [4:0] p5_bit_slice_13789_comb;
	wire [4:0] p5_concat_13790_comb;
	wire [4:0] p5_concat_13791_comb;
	wire [4:0] p5_concat_13792_comb;
	wire [4:0] p5_concat_13793_comb;
	wire [4:0] p5_bit_slice_13794_comb;
	wire [4:0] p5_concat_13795_comb;
	wire [4:0] p5_bit_slice_13796_comb;
	wire [4:0] p5_bit_slice_13797_comb;
	wire [4:0] p5_bit_slice_13798_comb;
	wire [4:0] p5_bit_slice_13799_comb;
	wire [4:0] p5_bit_slice_13800_comb;
	wire [4:0] p5_bit_slice_13801_comb;
	wire [4:0] p5_bit_slice_13802_comb;
	wire [4:0] p5_bit_slice_13803_comb;
	wire [21:0] p5_concat_13804_comb;
	wire [1:0] p5_bit_slice_13805_comb;
	wire [1:0] p5_bit_slice_13806_comb;
	wire [1:0] p5_bit_slice_13807_comb;
	wire [1:0] p5_bit_slice_13808_comb;
	wire [1:0] p5_bit_slice_13809_comb;
	wire [1:0] p5_bit_slice_13810_comb;
	wire [1:0] p5_bit_slice_13811_comb;
	wire [1:0] p5_concat_13812_comb;
	wire [1:0] p5_concat_13813_comb;
	wire [1:0] p5_concat_13814_comb;
	wire [1:0] p5_concat_13815_comb;
	wire [1:0] p5_bit_slice_13816_comb;
	wire [1:0] p5_bit_slice_13817_comb;
	wire [1:0] p5_concat_13818_comb;
	wire [1:0] p5_bit_slice_13819_comb;
	wire [1:0] p5_bit_slice_13820_comb;
	wire [1:0] p5_bit_slice_13821_comb;
	wire [1:0] p5_bit_slice_13822_comb;
	wire [1:0] p5_bit_slice_13823_comb;
	wire [1:0] p5_bit_slice_13824_comb;
	wire [1:0] p5_bit_slice_13825_comb;
	wire [20:0] p5_concat_13826_comb;
	wire p5_bit_slice_13827_comb;
	wire p5_bit_slice_13828_comb;
	wire p5_bit_slice_13829_comb;
	wire p5_bit_slice_13830_comb;
	wire p5_bit_slice_13831_comb;
	wire p5_bit_slice_13832_comb;
	wire p5_bit_slice_13833_comb;
	wire p5_bit_slice_13834_comb;
	wire p5_bit_slice_13835_comb;
	wire p5_bit_slice_13836_comb;
	wire p5_bit_slice_13837_comb;
	wire p5_bit_slice_13838_comb;
	wire p5_bit_slice_13839_comb;
	wire p5_bit_slice_13840_comb;
	wire p5_bit_slice_13841_comb;
	wire p5_bit_slice_13842_comb;
	wire p5_bit_slice_13843_comb;
	wire [5:0] p5_bit_slice_13844_comb;
	wire [5:0] p5_bit_slice_13845_comb;
	wire [5:0] p5_bit_slice_13846_comb;
	wire [5:0] p5_bit_slice_13847_comb;
	wire [5:0] p5_bit_slice_13848_comb;
	wire [5:0] p5_bit_slice_13849_comb;
	wire [5:0] p5_bit_slice_13850_comb;
	wire [5:0] p5_concat_13851_comb;
	wire [5:0] p5_bit_slice_13852_comb;
	wire [5:0] p5_concat_13853_comb;
	wire [5:0] p5_concat_13854_comb;
	wire [5:0] p5_bit_slice_13855_comb;
	wire [5:0] p5_concat_13856_comb;
	wire [5:0] p5_bit_slice_13857_comb;
	wire [5:0] p5_bit_slice_13858_comb;
	wire [5:0] p5_concat_13859_comb;
	wire [5:0] p5_bit_slice_13860_comb;
	wire [5:0] p5_bit_slice_13861_comb;
	wire [5:0] p5_bit_slice_13862_comb;
	wire [5:0] p5_concat_13863_comb;
	wire [5:0] p5_bit_slice_13864_comb;
	wire [5:0] p5_bit_slice_13865_comb;
	wire [21:0] p5_concat_13866_comb;
	wire [1:0] p5_bit_slice_13867_comb;
	wire [1:0] p5_bit_slice_13868_comb;
	wire [1:0] p5_bit_slice_13869_comb;
	wire [1:0] p5_bit_slice_13870_comb;
	wire [1:0] p5_bit_slice_13871_comb;
	wire [1:0] p5_bit_slice_13872_comb;
	wire [1:0] p5_concat_13873_comb;
	wire [1:0] p5_concat_13874_comb;
	wire [1:0] p5_concat_13875_comb;
	wire [1:0] p5_concat_13876_comb;
	wire [1:0] p5_concat_13877_comb;
	wire [1:0] p5_bit_slice_13878_comb;
	wire [1:0] p5_bit_slice_13879_comb;
	wire [1:0] p5_bit_slice_13880_comb;
	wire [1:0] p5_bit_slice_13881_comb;
	wire [1:0] p5_bit_slice_13882_comb;
	wire [1:0] p5_bit_slice_13883_comb;
	wire [1:0] p5_bit_slice_13884_comb;
	wire [1:0] p5_bit_slice_13885_comb;
	wire [1:0] p5_bit_slice_13886_comb;
	wire [1:0] p5_bit_slice_13887_comb;
	wire [1:0] p5_bit_slice_13888_comb;
	wire [22:0] p5_concat_13889_comb;
	wire [1:0] p5_bit_slice_13890_comb;
	wire [1:0] p5_bit_slice_13891_comb;
	wire [1:0] p5_bit_slice_13892_comb;
	wire [1:0] p5_bit_slice_13893_comb;
	wire [1:0] p5_bit_slice_13894_comb;
	wire [1:0] p5_bit_slice_13895_comb;
	wire [1:0] p5_bit_slice_13896_comb;
	wire [1:0] p5_bit_slice_13897_comb;
	wire [1:0] p5_concat_13898_comb;
	wire [1:0] p5_bit_slice_13899_comb;
	wire [1:0] p5_concat_13900_comb;
	wire [1:0] p5_concat_13901_comb;
	wire [1:0] p5_bit_slice_13902_comb;
	wire [1:0] p5_bit_slice_13903_comb;
	wire [1:0] p5_bit_slice_13904_comb;
	wire [1:0] p5_concat_13905_comb;
	wire [1:0] p5_bit_slice_13906_comb;
	wire [1:0] p5_bit_slice_13907_comb;
	wire [1:0] p5_bit_slice_13908_comb;
	wire [1:0] p5_bit_slice_13909_comb;
	wire [1:0] p5_xor_13910_comb;
	wire [1:0] p5_bit_slice_13911_comb;
	wire [1:0] p5_bit_slice_13912_comb;
	wire [21:0] p5_concat_13913_comb;
	wire [3:0] p5_bit_slice_13914_comb;
	wire [3:0] p5_bit_slice_13915_comb;
	wire [3:0] p5_bit_slice_13916_comb;
	wire [3:0] p5_bit_slice_13917_comb;
	wire [3:0] p5_bit_slice_13918_comb;
	wire [3:0] p5_bit_slice_13919_comb;
	wire [3:0] p5_bit_slice_13920_comb;
	wire [3:0] p5_bit_slice_13921_comb;
	wire [3:0] p5_concat_13922_comb;
	wire [3:0] p5_bit_slice_13923_comb;
	wire [3:0] p5_concat_13924_comb;
	wire [3:0] p5_concat_13925_comb;
	wire [3:0] p5_bit_slice_13926_comb;
	wire [3:0] p5_concat_13927_comb;
	wire [3:0] p5_bit_slice_13928_comb;
	wire [3:0] p5_bit_slice_13929_comb;
	wire [3:0] p5_bit_slice_13930_comb;
	wire [3:0] p5_bit_slice_13931_comb;
	wire [3:0] p5_bit_slice_13932_comb;
	wire [3:0] p5_bit_slice_13933_comb;
	wire [3:0] p5_bit_slice_13934_comb;
	wire [3:0] p5_bit_slice_13935_comb;
	wire [20:0] p5_concat_13936_comb;
	wire p5_bit_slice_13937_comb;
	wire p5_bit_slice_13938_comb;
	wire p5_bit_slice_13939_comb;
	wire p5_bit_slice_13940_comb;
	wire p5_bit_slice_13941_comb;
	wire p5_bit_slice_13942_comb;
	wire p5_bit_slice_13943_comb;
	wire p5_bit_slice_13944_comb;
	wire p5_bit_slice_13945_comb;
	wire p5_bit_slice_13946_comb;
	wire p5_bit_slice_13947_comb;
	wire p5_bit_slice_13948_comb;
	wire p5_bit_slice_13949_comb;
	wire p5_bit_slice_13950_comb;
	wire p5_bit_slice_13951_comb;
	wire p5_bit_slice_13952_comb;
	wire [20:0] p5_concat_13953_comb;
	wire [4:0] p5_bit_slice_13954_comb;
	wire [4:0] p5_bit_slice_13955_comb;
	wire [4:0] p5_bit_slice_13956_comb;
	wire [4:0] p5_bit_slice_13957_comb;
	wire [4:0] p5_bit_slice_13958_comb;
	wire [4:0] p5_bit_slice_13959_comb;
	wire [4:0] p5_bit_slice_13960_comb;
	wire [4:0] p5_concat_13961_comb;
	wire [4:0] p5_concat_13962_comb;
	wire [4:0] p5_concat_13963_comb;
	wire [4:0] p5_concat_13964_comb;
	wire [4:0] p5_bit_slice_13965_comb;
	wire [4:0] p5_bit_slice_13966_comb;
	wire [4:0] p5_bit_slice_13967_comb;
	wire [4:0] p5_concat_13968_comb;
	wire [4:0] p5_bit_slice_13969_comb;
	wire [4:0] p5_bit_slice_13970_comb;
	wire [4:0] p5_bit_slice_13971_comb;
	wire [4:0] p5_bit_slice_13972_comb;
	wire [4:0] p5_bit_slice_13973_comb;
	wire [21:0] p5_concat_13974_comb;
	wire [1:0] p5_bit_slice_13975_comb;
	wire [1:0] p5_bit_slice_13976_comb;
	wire [1:0] p5_bit_slice_13977_comb;
	wire [1:0] p5_bit_slice_13978_comb;
	wire [1:0] p5_bit_slice_13979_comb;
	wire [1:0] p5_bit_slice_13980_comb;
	wire [1:0] p5_bit_slice_13981_comb;
	wire [1:0] p5_concat_13982_comb;
	wire [1:0] p5_bit_slice_13983_comb;
	wire [1:0] p5_concat_13984_comb;
	wire [1:0] p5_concat_13985_comb;
	wire [1:0] p5_bit_slice_13986_comb;
	wire [1:0] p5_bit_slice_13987_comb;
	wire [1:0] p5_bit_slice_13988_comb;
	wire [1:0] p5_bit_slice_13989_comb;
	wire [1:0] p5_bit_slice_13990_comb;
	wire [1:0] p5_bit_slice_13991_comb;
	wire [1:0] p5_bit_slice_13992_comb;
	wire [1:0] p5_bit_slice_13993_comb;
	wire [1:0] p5_bit_slice_13994_comb;
	wire [1:0] p5_bit_slice_13995_comb;
	wire [1:0] p5_bit_slice_13996_comb;
	wire [19:0] p5_concat_13997_comb;
	wire p5_bit_slice_13998_comb;
	wire p5_bit_slice_13999_comb;
	wire p5_bit_slice_14000_comb;
	wire p5_bit_slice_14001_comb;
	wire p5_bit_slice_14002_comb;
	wire p5_bit_slice_14003_comb;
	wire p5_bit_slice_14004_comb;
	wire p5_bit_slice_14005_comb;
	wire p5_bit_slice_14006_comb;
	wire p5_bit_slice_14007_comb;
	wire p5_bit_slice_14008_comb;
	wire p5_bit_slice_14009_comb;
	wire p5_bit_slice_14010_comb;
	wire p5_bit_slice_14011_comb;
	wire p5_bit_slice_14012_comb;
	wire p5_bit_slice_14013_comb;
	wire p5_bit_slice_14014_comb;
	wire p5_one_hot_sel_14015_comb;
	wire [4:0] p5_one_hot_sel_14016_comb;
	wire [1:0] p5_one_hot_sel_14017_comb;
	wire p5_one_hot_sel_14018_comb;
	wire [5:0] p5_one_hot_sel_14019_comb;
	wire [1:0] p5_one_hot_sel_14020_comb;
	wire [1:0] p5_one_hot_sel_14021_comb;
	wire [3:0] p5_one_hot_sel_14022_comb;
	wire p5_one_hot_sel_14023_comb;
	wire [4:0] p5_one_hot_sel_14024_comb;
	wire [1:0] p5_one_hot_sel_14025_comb;
	wire p5_one_hot_sel_14026_comb;
	wire [31:0] p5_concat_14027_comb;
	wire [31:0] p5_sign_ext_14028_comb;
	wire [31:0] p5_and_14029_comb;
	wire [32:0] p5_tuple_14030_comb;
	assign p5_rotation_1__6_comb = p4_rs1[0];
	assign p5_rotation_1__5_comb = p4_rs1[31:1];
	assign p5_byte0__1_comb = p4_rs1[7:0];
	assign p5_rotation_2__5_comb = p4_rs1[31:8];
	assign p5_rotation_1__10_comb = p4_rs1[27:0];
	assign p5_rotation_1__9_comb = p4_rs1[31:28];
	assign p5_rotation_2__10_comb = p4_rs1[1:0];
	assign p5_rotation_2__9_comb = p4_rs1[31:2];
	assign p5_literal_13584_comb = 7'h00;
	assign p5_rotation_3__3_comb = p4_rs1[31:7];
	assign p5_rotation_1__1_comb = {p5_rotation_1__6_comb, p5_rotation_1__5_comb};
	assign p5_rotation_2__1_comb = {p5_byte0__1_comb, p5_rotation_2__5_comb};
	assign p5_rotation_1__2_comb = {p5_rotation_1__10_comb, p5_rotation_1__9_comb};
	assign p5_rotation_2__2_comb = {p5_rotation_2__10_comb, p5_rotation_2__9_comb};
	assign p5_rotation_3__4_comb = p4_rs1[6:0];
	assign p5_bit_slice_13591_comb = p4_rs1[27:26];
	assign p5_bit_slice_13592_comb = p4_rs1[6:5];
	assign p5_bit_slice_13593_comb = p4_rs1[25:21];
	assign p5_bit_slice_13594_comb = p4_rs1[31:27];
	assign p5_bit_slice_13595_comb = p4_rs1[4:0];
	assign p5_bit_slice_13596_comb = p4_rs1[12:11];
	assign p5_bit_slice_13597_comb = p4_rs1[21:20];
	assign p5_bit_slice_13598_comb = p4_rs1[31:21];
	assign p5_bit_slice_13599_comb = p4_rs1[10:0];
	assign p5_bit_slice_13600_comb = p4_rs1[19:9];
	assign p5_bit_slice_13601_comb = p4_rs1[6:4];
	assign p5_bit_slice_13602_comb = p4_rs1[17:15];
	assign p5_bit_slice_13603_comb = p4_rs1[3:0];
	assign p5_bit_slice_13604_comb = p4_rs1[14:11];
	assign p5_bit_slice_13605_comb = p4_rs1[20:0];
	assign p5_bit_slice_13606_comb = p4_rs1[26:6];
	assign p5_bit_slice_13607_comb = p4_rs1[31:11];
	assign p5_bit_slice_13608_comb = p4_rs1[27:17];
	assign p5_bit_slice_13609_comb = p4_rs1[20:12];
	assign p5_bit_slice_13610_comb = p4_rs1[31:23];
	assign p5_bit_slice_13611_comb = p4_rs1[8:0];
	assign p5_bit_slice_13612_comb = p4_rs1[18:14];
	assign p5_bit_slice_13613_comb = p4_rs1[26:13];
	assign p5_rotate_18__1_comb = p4_rs1[31:18];
	assign p5_bit_slice_13615_comb = p4_rs1[13:0];
	assign p5_bit_slice_13616_comb = p4_rs1[16:7];
	assign p5_bit_slice_13617_comb = p4_rs1[18:9];
	assign p5_bit_slice_13618_comb = p4_rs1[8:2];
	assign p5_rotation_3__5_comb = p4_rs1[31:25];
	assign p5_bit_slice_13620_comb = p4_rs1[20:7];
	assign p5_bit_slice_13621_comb = p4_rs1[16:3];
	assign p5_bit_slice_13622_comb = p4_rs1[11:2];
	assign p5_bit_slice_13623_comb = p4_rs1[22:13];
	assign p5_rot_c__1_comb = p4_rs1[31:22];
	assign p5_bit_slice_13625_comb = p4_rs1[5:2];
	assign p5_bit_slice_13626_comb = p4_rs1[10:7];
	assign p5_bit_slice_13627_comb = p4_rs1[12:6];
	assign p5_bit_slice_13628_comb = p4_rs1[17:11];
	assign p5_not_13629_comb = ~p4_rs1;
	assign p5_xor_13630_comb = p4_rs1 ^ p4_rs2;
	assign p5_shift_1_comb = {p5_literal_13584_comb, p5_rotation_3__3_comb};
	assign p5_combined_1_comb = p5_rotation_1__1_comb & p4_rs2;
	assign p5_combined_2_comb = p5_rotation_2__1_comb | p4_rs2;
	assign p5_rotation_1__12_comb = p4_rs1[5:0];
	assign p5_bit_slice_13635_comb = p4_rs1[10:5];
	assign p5_bit_slice_13636_comb = p4_rs1[24:19];
	assign p5_bit_slice_13637_comb = p4_rs1[28:23];
	assign p5_bit_slice_13638_comb = p4_rs2[18:13];
	assign p5_combined_1__1_comb = p5_rotation_1__2_comb & p4_rs2;
	assign p5_combined_2__1_comb = p5_rotation_2__2_comb | p4_rs2;
	assign p5_rotation_3__1_comb = {p5_rotation_3__4_comb, p5_rotation_3__3_comb};
	assign p5_bit_slice_13642_comb = p4_rs2[5:0];
	assign p5_bit_slice_13643_comb = p4_rs1[18:13];
	assign p5_or_13644_comb = p4_shll_13490 | p4_shrl_13491;
	assign p5_or_13645_comb = p4_shll_13492 | p4_shrl_13493;
	assign p5_result__44_comb = (p5_bit_slice_13591_comb ^ p5_rotation_2__10_comb) ^ p5_bit_slice_13592_comb;
	assign p5_result__43_comb = (p5_bit_slice_13593_comb ^ p5_bit_slice_13594_comb) ^ p5_bit_slice_13595_comb;
	assign p5_xor_13648_comb = (p5_rotation_2__10_comb ^ p5_bit_slice_13596_comb) ^ p5_bit_slice_13597_comb;
	assign p5_xor_13649_comb = (p5_bit_slice_13598_comb ^ p5_bit_slice_13599_comb) ^ p5_bit_slice_13600_comb;
	assign p5_xor_13650_comb = p5_bit_slice_13601_comb ^ p5_bit_slice_13602_comb;
	assign p5_xor_13651_comb = (p5_bit_slice_13603_comb ^ p5_bit_slice_13604_comb) ^ p5_rotation_1__9_comb;
	assign p5_result__42_comb = (p5_bit_slice_13605_comb ^ p5_bit_slice_13606_comb) ^ p5_bit_slice_13607_comb;
	assign p5_xor_13653_comb = (p5_bit_slice_13598_comb ^ p5_bit_slice_13599_comb) ^ p5_bit_slice_13608_comb;
	assign p5_bit_slice_13654_comb = p4_rs1[22:10];
	assign p5_rotation_1__13_comb = p4_rs1[31:19];
	assign p5_bit_slice_13656_comb = p4_rs2[12:0];
	assign p5_bit_slice_13657_comb = p4_rs1[12:0];
	assign p5_xor_13658_comb = (p5_bit_slice_13609_comb ^ p5_bit_slice_13610_comb) ^ p5_bit_slice_13611_comb;
	assign p5_xor_13659_comb = (p5_bit_slice_13594_comb ^ p5_bit_slice_13595_comb) ^ p5_bit_slice_13612_comb;
	assign p5_xor_13660_comb = (p5_bit_slice_13613_comb ^ p5_rotate_18__1_comb) ^ p5_bit_slice_13615_comb;
	assign p5_xor_13661_comb = p5_bit_slice_13616_comb ^ p5_bit_slice_13617_comb;
	assign p5_xor_13662_comb = (p5_rotation_3__4_comb ^ p5_bit_slice_13618_comb) ^ p5_rotation_3__5_comb;
	assign p5_xor_13663_comb = (p5_bit_slice_13620_comb ^ p5_rotate_18__1_comb) ^ p5_bit_slice_13621_comb;
	assign p5_xor_13664_comb = (p5_bit_slice_13622_comb ^ p5_bit_slice_13623_comb) ^ p5_rot_c__1_comb;
	assign p5_bit_slice_13665_comb = p4_rs1[9:0];
	assign p5_bit_slice_13666_comb = p4_rs1[29:17];
	assign p5_result__41_comb = (p5_rotation_1__9_comb ^ p5_bit_slice_13625_comb) ^ p5_bit_slice_13626_comb;
	assign p5_xor_13668_comb = (p5_bit_slice_13627_comb ^ p5_bit_slice_13628_comb) ^ p5_rotation_3__5_comb;
	assign p5_bit_slice_13669_comb = p4_rs1[8:6];
	assign p5_bit_slice_13670_comb = p4_rs1[21:19];
	assign p5_bit_slice_13671_comb = p4_rs2[31:29];
	assign p5_rotation_2__13_comb = p4_rs1[31:29];
	assign p5_or_13673_comb = p4_eq_13203 | p4_eq_13204;
	assign p5_or_13674_comb = p4_eq_13214 | p4_eq_13215;
	assign p5_or_13675_comb = p4_shrl_13494 | p4_shll_13495;
	assign p5_or_13676_comb = p4_shll_13496 | p4_shrl_13497;
	assign p5_or_13677_comb = p4_shrl_13498 | p4_shll_13499;
	assign p5_nor_13678_comb = ~(p5_not_13629_comb | p4_rs2);
	assign p5_nand_13679_comb = ~(p5_not_13629_comb & p4_rs2);
	assign p5_not_13680_comb = ~p5_xor_13630_comb;
	assign p5_xor_13681_comb = (((p5_rotation_1__1_comb ^ p5_rotation_2__1_comb) ^ p5_shift_1_comb) ^ p5_combined_1_comb) ^ p5_combined_2_comb;
	assign p5_xor_13682_comb = (p5_rotation_1__12_comb ^ p5_bit_slice_13635_comb) ^ p5_bit_slice_13636_comb;
	assign p5_xor_13683_comb = p5_bit_slice_13637_comb ^ p5_bit_slice_13638_comb;
	assign p5_xor_13684_comb = (((((p5_rotation_1__2_comb ^ p5_rotation_2__2_comb) ^ p5_rotation_3__1_comb) ^ p5_combined_1__1_comb) ^ p5_combined_2__1_comb) ^ p5_rotation_3__1_comb) ^ p4_rs2;
	assign p5_result__4_comb = (p5_bit_slice_13637_comb ^ p5_bit_slice_13642_comb) ^ p5_bit_slice_13638_comb;
	assign p5_xor_13686_comb = p5_bit_slice_13643_comb ^ p5_bit_slice_13637_comb;
	assign p5_result__7_comb = p4_rs1 ^ p5_or_13644_comb;
	assign p5_result__8_comb = p4_rs1 ^ p5_or_13645_comb;
	assign p5_result__28_comb = p4_rs1[25];
	assign p5_result__30_comb = p4_rs1[26];
	assign p5_result__32_comb = p4_rs1[27];
	assign p5_result__34_comb = p4_rs1[28];
	assign p5_result__36_comb = p4_rs1[29];
	assign p5_result__39_comb = p4_rs1[15];
	assign p5_result__38_comb = p4_rs1[30];
	assign p5_result__37_comb = p4_rs1[14];
	assign p5_result__35_comb = p4_rs1[13];
	assign p5_result__24_comb = p4_rs1[23];
	assign p5_result__20_comb = p4_rs1[21];
	assign p5_bit_slice_13700_comb = p5_result__44_comb[0];
	assign p5_bit_slice_13701_comb = p5_result__43_comb[4:1];
	assign p5_bit_slice_13702_comb = p5_xor_13648_comb[0];
	assign p5_bit_slice_13703_comb = p5_xor_13649_comb[10:7];
	assign p5_bit_slice_13704_comb = p5_xor_13650_comb[1:0];
	assign p5_bit_slice_13705_comb = p5_xor_13651_comb[3:1];
	assign p5_or_13706_comb = p4_eq_13223 | p4_eq_13224;
	assign p5_result__40_comb = p4_rs1[31];
	assign p5_result__33_comb = p4_rs1[12];
	assign p5_result__16_comb = p4_rs1[19];
	assign p5_result__12_comb = p4_rs1[17];
	assign p5_bit_slice_13711_comb = p5_result__43_comb[0];
	assign p5_bit_slice_13712_comb = p5_result__42_comb[20];
	assign p5_bit_slice_13713_comb = p5_xor_13651_comb[0];
	assign p5_bit_slice_13714_comb = p5_xor_13653_comb[10];
	assign p5_result__3_comb = (p5_bit_slice_13654_comb ^ p5_rotation_1__13_comb) ^ p5_bit_slice_13656_comb;
	assign p5_xor_13716_comb = (p5_bit_slice_13657_comb ^ p5_bit_slice_13654_comb) ^ p5_rotation_1__13_comb;
	assign p5_or_13717_comb = p4_eq_13225 | p4_eq_13215;
	assign p5_result__14_comb = p4_rs1[18];
	assign p5_result__18_comb = p4_rs1[20];
	assign p5_result__22_comb = p4_rs1[22];
	assign p5_result__31_comb = p4_rs1[11];
	assign p5_result__29_comb = p4_rs1[10];
	assign p5_result__27_comb = p4_rs1[9];
	assign p5_result__26_comb = p4_rs1[24];
	assign p5_result__23_comb = p4_rs1[7];
	assign p5_result__19_comb = p4_rs1[5];
	assign p5_result__15_comb = p4_rs1[3];
	assign p5_bit_slice_13728_comb = p5_xor_13649_comb[3:0];
	assign p5_bit_slice_13729_comb = p5_xor_13658_comb[8:7];
	assign p5_bit_slice_13730_comb = p5_xor_13659_comb[1:0];
	assign p5_bit_slice_13731_comb = p5_xor_13660_comb[13:10];
	assign p5_bit_slice_13732_comb = p5_xor_13661_comb[0];
	assign p5_bit_slice_13733_comb = p5_xor_13662_comb[6:2];
	assign p5_or_13734_comb = p4_eq_13225 | p4_eq_13214;
	assign p5_bit_slice_13735_comb = p4_rs2[0];
	assign p5_literal_13736_comb = 1'h0;
	assign p5_bit_slice_13737_comb = p4_rs2[7];
	assign p5_result__25_comb = p4_rs1[8];
	assign p5_result__11_comb = p4_rs1[1];
	assign p5_bit_slice_13740_comb = p5_xor_13653_comb[0];
	assign p5_bit_slice_13741_comb = p5_xor_13663_comb[13];
	assign p5_bit_slice_13742_comb = p4_rs1[31:30];
	assign p5_bit_slice_13743_comb = p4_rs1[24:23];
	assign p5_or_13744_comb = (p4_eq_13223 | p4_eq_13224) | p4_eq_13226;
	assign p5_result__21_comb = p4_rs1[6];
	assign p5_bit_slice_13746_comb = p5_xor_13658_comb[2:0];
	assign p5_bit_slice_13747_comb = p5_xor_13664_comb[9];
	assign p5_result__2_comb = (p5_bit_slice_13665_comb ^ p5_bit_slice_13617_comb) ^ p5_rot_c__1_comb;
	assign p5_xor_13749_comb = (p5_bit_slice_13666_comb ^ p5_rotation_1__13_comb) ^ p5_bit_slice_13654_comb;
	assign p5_result__13_comb = p4_rs1[2];
	assign p5_result__17_comb = p4_rs1[4];
	assign p5_bit_slice_13752_comb = p5_result__42_comb[3:0];
	assign p5_bit_slice_13753_comb = p5_result__41_comb[3];
	assign p5_bit_slice_13754_comb = p5_xor_13660_comb[0];
	assign p5_bit_slice_13755_comb = p5_xor_13668_comb[6:3];
	assign p5_result__10_comb = p4_rs1[16];
	assign p5_result__5_comb = (p5_bit_slice_13669_comb ^ p5_bit_slice_13670_comb) ^ p5_bit_slice_13671_comb;
	assign p5_xor_13758_comb = (p5_bit_slice_13670_comb ^ p5_rotation_2__13_comb) ^ p5_bit_slice_13669_comb;
	assign p5_or_13759_comb = (p5_or_13673_comb | p4_eq_13214) | p4_eq_13215;
	assign p5_concat_13760_comb = {p4_eq_13227, p4_eq_13228, p4_eq_13229, p4_eq_13226, p4_eq_13224, p4_eq_13230, p4_eq_13223, p4_eq_13231, p4_eq_13232, p4_eq_13233, p4_eq_13234, p4_eq_13235, p5_or_13674_comb, p4_eq_13225, p4_eq_13236, p4_eq_13203, p4_eq_13237, p4_eq_13238, p4_eq_13239, p4_eq_13240, p4_eq_13241, p4_eq_13242};
	assign p5_bit_slice_13761_comb = p5_or_13675_comb[31];
	assign p5_bit_slice_13762_comb = p5_or_13676_comb[31];
	assign p5_bit_slice_13763_comb = p5_or_13677_comb[31];
	assign p5_bit_slice_13764_comb = p5_nor_13678_comb[31];
	assign p5_bit_slice_13765_comb = p5_nand_13679_comb[31];
	assign p5_bit_slice_13766_comb = p5_not_13680_comb[31];
	assign p5_bit_slice_13767_comb = p4_rs2[15];
	assign p5_bit_slice_13768_comb = p5_result__44_comb[1];
	assign p5_bit_slice_13769_comb = p5_xor_13648_comb[1];
	assign p5_bit_slice_13770_comb = p5_xor_13681_comb[31];
	assign p5_bit_slice_13771_comb = p5_xor_13650_comb[2];
	assign p5_bit_slice_13772_comb = p5_xor_13682_comb[5];
	assign p5_bit_slice_13773_comb = p5_xor_13683_comb[5];
	assign p5_bit_slice_13774_comb = p5_xor_13684_comb[31];
	assign p5_bit_slice_13775_comb = p5_result__4_comb[5];
	assign p5_bit_slice_13776_comb = p5_xor_13686_comb[5];
	assign p5_bit_slice_13777_comb = p5_xor_13661_comb[9];
	assign p5_bit_slice_13778_comb = p5_result__7_comb[31];
	assign p5_bit_slice_13779_comb = p5_result__8_comb[31];
	assign p5_concat_13780_comb = {p4_eq_13227, p4_eq_13228, p4_eq_13229, p4_eq_13226, p4_eq_13224, p4_eq_13230, p4_eq_13223, p4_eq_13231, p4_eq_13232, p4_eq_13233, p4_eq_13234, p4_eq_13235, p4_eq_13215, p4_eq_13214, p4_eq_13225, p4_eq_13236, p4_eq_13203, p4_eq_13237, p4_eq_13238, p4_eq_13239, p4_eq_13240, p4_eq_13241, p4_eq_13242};
	assign p5_bit_slice_13781_comb = p5_or_13675_comb[30:26];
	assign p5_bit_slice_13782_comb = p5_or_13676_comb[30:26];
	assign p5_bit_slice_13783_comb = p5_or_13677_comb[30:26];
	assign p5_bit_slice_13784_comb = p5_nor_13678_comb[30:26];
	assign p5_bit_slice_13785_comb = p5_nand_13679_comb[30:26];
	assign p5_bit_slice_13786_comb = p5_not_13680_comb[30:26];
	assign p5_bit_slice_13787_comb = p4_rs2[14:10];
	assign p5_concat_13788_comb = {p5_result__28_comb, p5_result__30_comb, p5_result__32_comb, p5_result__34_comb, p5_result__36_comb};
	assign p5_bit_slice_13789_comb = p4_rs1[6:2];
	assign p5_concat_13790_comb = {p5_result__39_comb, p5_result__38_comb, p5_result__37_comb, p5_result__36_comb, p5_result__35_comb};
	assign p5_concat_13791_comb = {p5_result__36_comb, p5_result__32_comb, p5_result__28_comb, p5_result__24_comb, p5_result__20_comb};
	assign p5_concat_13792_comb = {p5_bit_slice_13700_comb, p5_bit_slice_13701_comb};
	assign p5_concat_13793_comb = {p5_bit_slice_13702_comb, p5_bit_slice_13703_comb};
	assign p5_bit_slice_13794_comb = p5_xor_13681_comb[30:26];
	assign p5_concat_13795_comb = {p5_bit_slice_13704_comb, p5_bit_slice_13705_comb};
	assign p5_bit_slice_13796_comb = p5_xor_13682_comb[4:0];
	assign p5_bit_slice_13797_comb = p5_xor_13683_comb[4:0];
	assign p5_bit_slice_13798_comb = p5_xor_13684_comb[30:26];
	assign p5_bit_slice_13799_comb = p5_result__4_comb[4:0];
	assign p5_bit_slice_13800_comb = p5_xor_13686_comb[4:0];
	assign p5_bit_slice_13801_comb = p5_xor_13661_comb[8:4];
	assign p5_bit_slice_13802_comb = p5_result__7_comb[30:26];
	assign p5_bit_slice_13803_comb = p5_result__8_comb[30:26];
	assign p5_concat_13804_comb = {p4_eq_13227, p4_eq_13228, p4_eq_13229, p4_eq_13226, p4_eq_13230, p5_or_13706_comb, p4_eq_13231, p4_eq_13232, p4_eq_13233, p4_eq_13234, p4_eq_13235, p4_eq_13215, p4_eq_13214, p4_eq_13225, p4_eq_13236, p4_eq_13203, p4_eq_13237, p4_eq_13238, p4_eq_13239, p4_eq_13240, p4_eq_13241, p4_eq_13242};
	assign p5_bit_slice_13805_comb = p5_or_13675_comb[25:24];
	assign p5_bit_slice_13806_comb = p5_or_13676_comb[25:24];
	assign p5_bit_slice_13807_comb = p5_or_13677_comb[25:24];
	assign p5_bit_slice_13808_comb = p5_nor_13678_comb[25:24];
	assign p5_bit_slice_13809_comb = p5_nand_13679_comb[25:24];
	assign p5_bit_slice_13810_comb = p5_not_13680_comb[25:24];
	assign p5_bit_slice_13811_comb = p4_rs2[9:8];
	assign p5_concat_13812_comb = {p5_result__38_comb, p5_result__40_comb};
	assign p5_concat_13813_comb = {p5_result__34_comb, p5_result__33_comb};
	assign p5_concat_13814_comb = {p5_result__16_comb, p5_result__12_comb};
	assign p5_concat_13815_comb = {p5_bit_slice_13711_comb, p5_bit_slice_13712_comb};
	assign p5_bit_slice_13816_comb = p5_xor_13649_comb[6:5];
	assign p5_bit_slice_13817_comb = p5_xor_13681_comb[25:24];
	assign p5_concat_13818_comb = {p5_bit_slice_13713_comb, p5_bit_slice_13714_comb};
	assign p5_bit_slice_13819_comb = p5_xor_13659_comb[4:3];
	assign p5_bit_slice_13820_comb = p5_result__3_comb[12:11];
	assign p5_bit_slice_13821_comb = p5_xor_13684_comb[25:24];
	assign p5_bit_slice_13822_comb = p5_xor_13716_comb[12:11];
	assign p5_bit_slice_13823_comb = p5_xor_13661_comb[3:2];
	assign p5_bit_slice_13824_comb = p5_result__7_comb[25:24];
	assign p5_bit_slice_13825_comb = p5_result__8_comb[25:24];
	assign p5_concat_13826_comb = {p4_eq_13227, p4_eq_13228, p4_eq_13229, p4_eq_13226, p4_eq_13230, p5_or_13706_comb, p4_eq_13231, p4_eq_13232, p4_eq_13233, p4_eq_13234, p4_eq_13235, p4_eq_13214, p5_or_13717_comb, p4_eq_13236, p4_eq_13203, p4_eq_13237, p4_eq_13238, p4_eq_13239, p4_eq_13240, p4_eq_13241, p4_eq_13242};
	assign p5_bit_slice_13827_comb = p5_or_13675_comb[23];
	assign p5_bit_slice_13828_comb = p5_or_13676_comb[23];
	assign p5_bit_slice_13829_comb = p5_or_13677_comb[23];
	assign p5_bit_slice_13830_comb = p5_nor_13678_comb[23];
	assign p5_bit_slice_13831_comb = p5_nand_13679_comb[23];
	assign p5_bit_slice_13832_comb = p5_not_13680_comb[23];
	assign p5_bit_slice_13833_comb = p5_result__42_comb[19];
	assign p5_bit_slice_13834_comb = p5_xor_13649_comb[4];
	assign p5_bit_slice_13835_comb = p5_xor_13681_comb[23];
	assign p5_bit_slice_13836_comb = p5_xor_13653_comb[9];
	assign p5_bit_slice_13837_comb = p5_xor_13659_comb[2];
	assign p5_bit_slice_13838_comb = p5_result__3_comb[10];
	assign p5_bit_slice_13839_comb = p5_xor_13684_comb[23];
	assign p5_bit_slice_13840_comb = p5_xor_13716_comb[10];
	assign p5_bit_slice_13841_comb = p5_xor_13661_comb[1];
	assign p5_bit_slice_13842_comb = p5_result__7_comb[23];
	assign p5_bit_slice_13843_comb = p5_result__8_comb[23];
	assign p5_bit_slice_13844_comb = p5_or_13675_comb[22:17];
	assign p5_bit_slice_13845_comb = p5_or_13676_comb[22:17];
	assign p5_bit_slice_13846_comb = p5_or_13677_comb[22:17];
	assign p5_bit_slice_13847_comb = p5_nor_13678_comb[22:17];
	assign p5_bit_slice_13848_comb = p5_nand_13679_comb[22:17];
	assign p5_bit_slice_13849_comb = p5_not_13680_comb[22:17];
	assign p5_bit_slice_13850_comb = p4_rs2[6:1];
	assign p5_concat_13851_comb = {p5_result__12_comb, p5_result__14_comb, p5_result__16_comb, p5_result__18_comb, p5_result__20_comb, p5_result__22_comb};
	assign p5_bit_slice_13852_comb = p4_rs1[14:9];
	assign p5_concat_13853_comb = {p5_result__31_comb, p5_result__30_comb, p5_result__29_comb, p5_result__28_comb, p5_result__27_comb, p5_result__26_comb};
	assign p5_concat_13854_comb = {p5_result__35_comb, p5_result__31_comb, p5_result__27_comb, p5_result__23_comb, p5_result__19_comb, p5_result__15_comb};
	assign p5_bit_slice_13855_comb = p5_result__42_comb[18:13];
	assign p5_concat_13856_comb = {p5_bit_slice_13728_comb, p5_bit_slice_13729_comb};
	assign p5_bit_slice_13857_comb = p5_xor_13681_comb[22:17];
	assign p5_bit_slice_13858_comb = p5_xor_13653_comb[8:3];
	assign p5_concat_13859_comb = {p5_bit_slice_13730_comb, p5_bit_slice_13731_comb};
	assign p5_bit_slice_13860_comb = p5_result__3_comb[9:4];
	assign p5_bit_slice_13861_comb = p5_xor_13684_comb[22:17];
	assign p5_bit_slice_13862_comb = p5_xor_13716_comb[9:4];
	assign p5_concat_13863_comb = {p5_bit_slice_13732_comb, p5_bit_slice_13733_comb};
	assign p5_bit_slice_13864_comb = p5_result__7_comb[22:17];
	assign p5_bit_slice_13865_comb = p5_result__8_comb[22:17];
	assign p5_concat_13866_comb = {p4_eq_13227, p4_eq_13228, p4_eq_13229, p4_eq_13226, p4_eq_13230, p5_or_13706_comb, p4_eq_13231, p4_eq_13232, p4_eq_13233, p4_eq_13234, p4_eq_13235, p4_eq_13215, p5_or_13734_comb, p4_eq_13236, p4_eq_13204, p4_eq_13203, p4_eq_13237, p4_eq_13238, p4_eq_13239, p4_eq_13240, p4_eq_13241, p4_eq_13242};
	assign p5_bit_slice_13867_comb = p5_or_13675_comb[16:15];
	assign p5_bit_slice_13868_comb = p5_or_13676_comb[16:15];
	assign p5_bit_slice_13869_comb = p5_or_13677_comb[16:15];
	assign p5_bit_slice_13870_comb = p5_nor_13678_comb[16:15];
	assign p5_bit_slice_13871_comb = p5_nand_13679_comb[16:15];
	assign p5_bit_slice_13872_comb = p5_not_13680_comb[16:15];
	assign p5_concat_13873_comb = {p5_bit_slice_13735_comb, p5_result__39_comb};
	assign p5_concat_13874_comb = {p5_literal_13736_comb, p5_bit_slice_13737_comb};
	assign p5_concat_13875_comb = {p5_result__24_comb, p5_result__25_comb};
	assign p5_concat_13876_comb = {p5_result__25_comb, p5_result__24_comb};
	assign p5_concat_13877_comb = {p5_result__11_comb, p5_result__38_comb};
	assign p5_bit_slice_13878_comb = p5_result__42_comb[12:11];
	assign p5_bit_slice_13879_comb = p5_xor_13658_comb[6:5];
	assign p5_bit_slice_13880_comb = p5_xor_13681_comb[16:15];
	assign p5_bit_slice_13881_comb = p5_xor_13653_comb[2:1];
	assign p5_bit_slice_13882_comb = p5_xor_13660_comb[9:8];
	assign p5_bit_slice_13883_comb = p5_result__3_comb[3:2];
	assign p5_bit_slice_13884_comb = p5_xor_13684_comb[16:15];
	assign p5_bit_slice_13885_comb = p5_xor_13716_comb[3:2];
	assign p5_bit_slice_13886_comb = p5_xor_13662_comb[1:0];
	assign p5_bit_slice_13887_comb = p5_result__7_comb[16:15];
	assign p5_bit_slice_13888_comb = p5_result__8_comb[16:15];
	assign p5_concat_13889_comb = {p4_eq_13227, p4_eq_13228, p4_eq_13229, p4_eq_13226, p4_eq_13230, p5_or_13706_comb, p4_eq_13231, p4_eq_13232, p4_eq_13233, p4_eq_13234, p4_eq_13235, p4_eq_13215, p4_eq_13214, p4_eq_13225, p4_eq_13236, p4_eq_13204, p4_eq_13203, p4_eq_13237, p4_eq_13238, p4_eq_13239, p4_eq_13240, p4_eq_13241, p4_eq_13242};
	assign p5_bit_slice_13890_comb = p5_or_13675_comb[14:13];
	assign p5_bit_slice_13891_comb = p5_or_13676_comb[14:13];
	assign p5_bit_slice_13892_comb = p5_or_13677_comb[14:13];
	assign p5_bit_slice_13893_comb = p5_nor_13678_comb[14:13];
	assign p5_bit_slice_13894_comb = p5_nand_13679_comb[14:13];
	assign p5_bit_slice_13895_comb = p5_not_13680_comb[14:13];
	assign p5_bit_slice_13896_comb = p4_rs1[14:13];
	assign p5_bit_slice_13897_comb = p4_rs2[6:5];
	assign p5_concat_13898_comb = {p5_result__27_comb, p5_result__29_comb};
	assign p5_bit_slice_13899_comb = p4_rs1[22:21];
	assign p5_concat_13900_comb = {p5_result__23_comb, p5_result__22_comb};
	assign p5_concat_13901_comb = {p5_result__34_comb, p5_result__30_comb};
	assign p5_bit_slice_13902_comb = p5_result__42_comb[10:9];
	assign p5_bit_slice_13903_comb = p5_xor_13658_comb[4:3];
	assign p5_bit_slice_13904_comb = p5_xor_13681_comb[14:13];
	assign p5_concat_13905_comb = {p5_bit_slice_13740_comb, p5_bit_slice_13741_comb};
	assign p5_bit_slice_13906_comb = p5_xor_13660_comb[7:6];
	assign p5_bit_slice_13907_comb = p5_result__3_comb[1:0];
	assign p5_bit_slice_13908_comb = p5_xor_13684_comb[14:13];
	assign p5_bit_slice_13909_comb = p5_xor_13716_comb[1:0];
	assign p5_xor_13910_comb = (p5_bit_slice_13742_comb ^ p5_rotation_2__10_comb) ^ p5_bit_slice_13743_comb;
	assign p5_bit_slice_13911_comb = p5_result__7_comb[14:13];
	assign p5_bit_slice_13912_comb = p5_result__8_comb[14:13];
	assign p5_concat_13913_comb = {p4_eq_13227, p4_eq_13228, p4_eq_13229, p4_eq_13230, p5_or_13744_comb, p4_eq_13231, p4_eq_13232, p4_eq_13233, p4_eq_13234, p4_eq_13235, p4_eq_13215, p4_eq_13214, p4_eq_13225, p4_eq_13236, p4_eq_13204, p4_eq_13203, p4_eq_13237, p4_eq_13238, p4_eq_13239, p4_eq_13240, p4_eq_13241, p4_eq_13242};
	assign p5_bit_slice_13914_comb = p5_or_13675_comb[12:9];
	assign p5_bit_slice_13915_comb = p5_or_13676_comb[12:9];
	assign p5_bit_slice_13916_comb = p5_or_13677_comb[12:9];
	assign p5_bit_slice_13917_comb = p5_nor_13678_comb[12:9];
	assign p5_bit_slice_13918_comb = p5_nand_13679_comb[12:9];
	assign p5_bit_slice_13919_comb = p5_not_13680_comb[12:9];
	assign p5_bit_slice_13920_comb = p4_rs1[12:9];
	assign p5_bit_slice_13921_comb = p4_rs2[4:1];
	assign p5_concat_13922_comb = {p5_result__31_comb, p5_result__33_comb, p5_result__35_comb, p5_result__37_comb};
	assign p5_bit_slice_13923_comb = p4_rs1[20:17];
	assign p5_concat_13924_comb = {p5_result__21_comb, p5_result__20_comb, p5_result__19_comb, p5_result__18_comb};
	assign p5_concat_13925_comb = {p5_result__26_comb, p5_result__22_comb, p5_result__18_comb, p5_result__14_comb};
	assign p5_bit_slice_13926_comb = p5_result__42_comb[8:5];
	assign p5_concat_13927_comb = {p5_bit_slice_13746_comb, p5_bit_slice_13747_comb};
	assign p5_bit_slice_13928_comb = p5_xor_13681_comb[12:9];
	assign p5_bit_slice_13929_comb = p5_xor_13663_comb[12:9];
	assign p5_bit_slice_13930_comb = p5_xor_13660_comb[5:2];
	assign p5_bit_slice_13931_comb = p5_result__2_comb[9:6];
	assign p5_bit_slice_13932_comb = p5_xor_13684_comb[12:9];
	assign p5_bit_slice_13933_comb = p5_xor_13749_comb[12:9];
	assign p5_bit_slice_13934_comb = p5_result__7_comb[12:9];
	assign p5_bit_slice_13935_comb = p5_result__8_comb[12:9];
	assign p5_concat_13936_comb = {p4_eq_13227, p4_eq_13228, p4_eq_13229, p4_eq_13230, p5_or_13744_comb, p4_eq_13231, p4_eq_13232, p4_eq_13233, p4_eq_13234, p4_eq_13235, p4_eq_13214, p5_or_13717_comb, p4_eq_13236, p4_eq_13204, p4_eq_13203, p4_eq_13237, p4_eq_13238, p4_eq_13239, p4_eq_13240, p4_eq_13241, p4_eq_13242};
	assign p5_bit_slice_13937_comb = p5_or_13675_comb[8];
	assign p5_bit_slice_13938_comb = p5_or_13676_comb[8];
	assign p5_bit_slice_13939_comb = p5_or_13677_comb[8];
	assign p5_bit_slice_13940_comb = p5_nor_13678_comb[8];
	assign p5_bit_slice_13941_comb = p5_nand_13679_comb[8];
	assign p5_bit_slice_13942_comb = p5_not_13680_comb[8];
	assign p5_bit_slice_13943_comb = p5_result__42_comb[4];
	assign p5_bit_slice_13944_comb = p5_xor_13664_comb[8];
	assign p5_bit_slice_13945_comb = p5_xor_13681_comb[8];
	assign p5_bit_slice_13946_comb = p5_xor_13663_comb[8];
	assign p5_bit_slice_13947_comb = p5_xor_13660_comb[1];
	assign p5_bit_slice_13948_comb = p5_result__2_comb[5];
	assign p5_bit_slice_13949_comb = p5_xor_13684_comb[8];
	assign p5_bit_slice_13950_comb = p5_xor_13749_comb[8];
	assign p5_bit_slice_13951_comb = p5_result__7_comb[8];
	assign p5_bit_slice_13952_comb = p5_result__8_comb[8];
	assign p5_concat_13953_comb = {p4_eq_13227, p4_eq_13228, p4_eq_13229, p4_eq_13230, p5_or_13744_comb, p4_eq_13231, p4_eq_13232, p4_eq_13233, p4_eq_13234, p4_eq_13235, p4_eq_13215, p4_eq_13214, p4_eq_13225, p4_eq_13236, p5_or_13673_comb, p4_eq_13237, p4_eq_13238, p4_eq_13239, p4_eq_13240, p4_eq_13241, p4_eq_13242};
	assign p5_bit_slice_13954_comb = p5_or_13675_comb[7:3];
	assign p5_bit_slice_13955_comb = p5_or_13676_comb[7:3];
	assign p5_bit_slice_13956_comb = p5_or_13677_comb[7:3];
	assign p5_bit_slice_13957_comb = p5_nor_13678_comb[7:3];
	assign p5_bit_slice_13958_comb = p5_nand_13679_comb[7:3];
	assign p5_bit_slice_13959_comb = p5_not_13680_comb[7:3];
	assign p5_bit_slice_13960_comb = p4_rs1[7:3];
	assign p5_concat_13961_comb = {p5_rotation_1__6_comb, p5_result__11_comb, p5_result__13_comb, p5_result__15_comb, p5_result__17_comb};
	assign p5_concat_13962_comb = {p5_result__16_comb, p5_result__15_comb, p5_result__14_comb, p5_result__13_comb, p5_result__12_comb};
	assign p5_concat_13963_comb = {p5_result__37_comb, p5_result__33_comb, p5_result__29_comb, p5_result__25_comb, p5_result__21_comb};
	assign p5_concat_13964_comb = {p5_bit_slice_13752_comb, p5_bit_slice_13753_comb};
	assign p5_bit_slice_13965_comb = p5_xor_13664_comb[7:3];
	assign p5_bit_slice_13966_comb = p5_xor_13681_comb[7:3];
	assign p5_bit_slice_13967_comb = p5_xor_13663_comb[7:3];
	assign p5_concat_13968_comb = {p5_bit_slice_13754_comb, p5_bit_slice_13755_comb};
	assign p5_bit_slice_13969_comb = p5_result__2_comb[4:0];
	assign p5_bit_slice_13970_comb = p5_xor_13684_comb[7:3];
	assign p5_bit_slice_13971_comb = p5_xor_13749_comb[7:3];
	assign p5_bit_slice_13972_comb = p5_result__7_comb[7:3];
	assign p5_bit_slice_13973_comb = p5_result__8_comb[7:3];
	assign p5_concat_13974_comb = {p4_eq_13227, p4_eq_13228, p4_eq_13229, p4_eq_13226, p4_eq_13230, p5_or_13706_comb, p4_eq_13231, p4_eq_13232, p4_eq_13233, p4_eq_13234, p4_eq_13235, p4_eq_13215, p4_eq_13214, p4_eq_13225, p4_eq_13236, p5_or_13673_comb, p4_eq_13237, p4_eq_13238, p4_eq_13239, p4_eq_13240, p4_eq_13241, p4_eq_13242};
	assign p5_bit_slice_13975_comb = p5_or_13675_comb[2:1];
	assign p5_bit_slice_13976_comb = p5_or_13676_comb[2:1];
	assign p5_bit_slice_13977_comb = p5_or_13677_comb[2:1];
	assign p5_bit_slice_13978_comb = p5_nor_13678_comb[2:1];
	assign p5_bit_slice_13979_comb = p5_nand_13679_comb[2:1];
	assign p5_bit_slice_13980_comb = p5_not_13680_comb[2:1];
	assign p5_bit_slice_13981_comb = p4_rs1[2:1];
	assign p5_concat_13982_comb = {p5_result__19_comb, p5_result__21_comb};
	assign p5_bit_slice_13983_comb = p4_rs1[26:25];
	assign p5_concat_13984_comb = {p5_result__11_comb, p5_result__10_comb};
	assign p5_concat_13985_comb = {p5_result__17_comb, p5_result__13_comb};
	assign p5_bit_slice_13986_comb = p5_result__41_comb[2:1];
	assign p5_bit_slice_13987_comb = p5_xor_13664_comb[2:1];
	assign p5_bit_slice_13988_comb = p5_xor_13681_comb[2:1];
	assign p5_bit_slice_13989_comb = p5_xor_13663_comb[2:1];
	assign p5_bit_slice_13990_comb = p5_xor_13668_comb[2:1];
	assign p5_bit_slice_13991_comb = p5_result__5_comb[2:1];
	assign p5_bit_slice_13992_comb = p5_xor_13684_comb[2:1];
	assign p5_bit_slice_13993_comb = p5_xor_13758_comb[2:1];
	assign p5_bit_slice_13994_comb = p5_xor_13749_comb[2:1];
	assign p5_bit_slice_13995_comb = p5_result__7_comb[2:1];
	assign p5_bit_slice_13996_comb = p5_result__8_comb[2:1];
	assign p5_concat_13997_comb = {p4_eq_13227, p4_eq_13228, p4_eq_13229, p4_eq_13226, p4_eq_13230, p5_or_13706_comb, p4_eq_13231, p4_eq_13232, p4_eq_13233, p4_eq_13234, p4_eq_13235, p4_eq_13225, p4_eq_13236, p5_or_13759_comb, p4_eq_13237, p4_eq_13238, p4_eq_13239, p4_eq_13240, p4_eq_13241, p4_eq_13242};
	assign p5_bit_slice_13998_comb = p5_or_13675_comb[0];
	assign p5_bit_slice_13999_comb = p5_or_13676_comb[0];
	assign p5_bit_slice_14000_comb = p5_or_13677_comb[0];
	assign p5_bit_slice_14001_comb = p5_nor_13678_comb[0];
	assign p5_bit_slice_14002_comb = p5_nand_13679_comb[0];
	assign p5_bit_slice_14003_comb = p5_not_13680_comb[0];
	assign p5_bit_slice_14004_comb = p5_result__41_comb[0];
	assign p5_bit_slice_14005_comb = p5_xor_13664_comb[0];
	assign p5_bit_slice_14006_comb = p5_xor_13681_comb[0];
	assign p5_bit_slice_14007_comb = p5_xor_13663_comb[0];
	assign p5_bit_slice_14008_comb = p5_xor_13668_comb[0];
	assign p5_bit_slice_14009_comb = p5_result__5_comb[0];
	assign p5_bit_slice_14010_comb = p5_xor_13684_comb[0];
	assign p5_bit_slice_14011_comb = p5_xor_13758_comb[0];
	assign p5_bit_slice_14012_comb = p5_xor_13749_comb[0];
	assign p5_bit_slice_14013_comb = p5_result__7_comb[0];
	assign p5_bit_slice_14014_comb = p5_result__8_comb[0];
	assign p5_one_hot_sel_14015_comb = (((((((((((((((((((((p5_bit_slice_13761_comb & p5_concat_13760_comb[0]) | (p5_bit_slice_13762_comb & p5_concat_13760_comb[1])) | (p5_bit_slice_13763_comb & p5_concat_13760_comb[2])) | (p5_bit_slice_13764_comb & p5_concat_13760_comb[3])) | (p5_bit_slice_13765_comb & p5_concat_13760_comb[4])) | (p5_bit_slice_13766_comb & p5_concat_13760_comb[5])) | (p5_bit_slice_13767_comb & p5_concat_13760_comb[6])) | (p5_result__26_comb & p5_concat_13760_comb[7])) | (p5_result__23_comb & p5_concat_13760_comb[8])) | (p5_result__40_comb & p5_concat_13760_comb[9])) | (p5_bit_slice_13768_comb & p5_concat_13760_comb[10])) | (p5_bit_slice_13769_comb & p5_concat_13760_comb[11])) | (p5_bit_slice_13770_comb & p5_concat_13760_comb[12])) | (p5_bit_slice_13771_comb & p5_concat_13760_comb[13])) | (p5_bit_slice_13772_comb & p5_concat_13760_comb[14])) | (p5_bit_slice_13773_comb & p5_concat_13760_comb[15])) | (p5_bit_slice_13774_comb & p5_concat_13760_comb[16])) | (p5_bit_slice_13775_comb & p5_concat_13760_comb[17])) | (p5_bit_slice_13776_comb & p5_concat_13760_comb[18])) | (p5_bit_slice_13777_comb & p5_concat_13760_comb[19])) | (p5_bit_slice_13778_comb & p5_concat_13760_comb[20])) | (p5_bit_slice_13779_comb & p5_concat_13760_comb[21]);
	assign p5_one_hot_sel_14016_comb = ((((((((((((((((((((((p5_bit_slice_13781_comb & {5 {p5_concat_13780_comb[0]}}) | (p5_bit_slice_13782_comb & {5 {p5_concat_13780_comb[1]}})) | (p5_bit_slice_13783_comb & {5 {p5_concat_13780_comb[2]}})) | (p5_bit_slice_13784_comb & {5 {p5_concat_13780_comb[3]}})) | (p5_bit_slice_13785_comb & {5 {p5_concat_13780_comb[4]}})) | (p5_bit_slice_13786_comb & {5 {p5_concat_13780_comb[5]}})) | (p5_bit_slice_13787_comb & {5 {p5_concat_13780_comb[6]}})) | (p5_concat_13788_comb & {5 {p5_concat_13780_comb[7]}})) | (p5_bit_slice_13789_comb & {5 {p5_concat_13780_comb[8]}})) | (p5_concat_13790_comb & {5 {p5_concat_13780_comb[9]}})) | (p5_concat_13791_comb & {5 {p5_concat_13780_comb[10]}})) | (p5_concat_13792_comb & {5 {p5_concat_13780_comb[11]}})) | (p5_concat_13793_comb & {5 {p5_concat_13780_comb[12]}})) | (p5_bit_slice_13794_comb & {5 {p5_concat_13780_comb[13]}})) | (p5_concat_13795_comb & {5 {p5_concat_13780_comb[14]}})) | (p5_bit_slice_13796_comb & {5 {p5_concat_13780_comb[15]}})) | (p5_bit_slice_13797_comb & {5 {p5_concat_13780_comb[16]}})) | (p5_bit_slice_13798_comb & {5 {p5_concat_13780_comb[17]}})) | (p5_bit_slice_13799_comb & {5 {p5_concat_13780_comb[18]}})) | (p5_bit_slice_13800_comb & {5 {p5_concat_13780_comb[19]}})) | (p5_bit_slice_13801_comb & {5 {p5_concat_13780_comb[20]}})) | (p5_bit_slice_13802_comb & {5 {p5_concat_13780_comb[21]}})) | (p5_bit_slice_13803_comb & {5 {p5_concat_13780_comb[22]}});
	assign p5_one_hot_sel_14017_comb = (((((((((((((((((((((p5_bit_slice_13805_comb & {2 {p5_concat_13804_comb[0]}}) | (p5_bit_slice_13806_comb & {2 {p5_concat_13804_comb[1]}})) | (p5_bit_slice_13807_comb & {2 {p5_concat_13804_comb[2]}})) | (p5_bit_slice_13808_comb & {2 {p5_concat_13804_comb[3]}})) | (p5_bit_slice_13809_comb & {2 {p5_concat_13804_comb[4]}})) | (p5_bit_slice_13810_comb & {2 {p5_concat_13804_comb[5]}})) | (p5_bit_slice_13811_comb & {2 {p5_concat_13804_comb[6]}})) | (p5_concat_13812_comb & {2 {p5_concat_13804_comb[7]}})) | (p5_rotation_2__10_comb & {2 {p5_concat_13804_comb[8]}})) | (p5_concat_13813_comb & {2 {p5_concat_13804_comb[9]}})) | (p5_concat_13814_comb & {2 {p5_concat_13804_comb[10]}})) | (p5_concat_13815_comb & {2 {p5_concat_13804_comb[11]}})) | (p5_bit_slice_13816_comb & {2 {p5_concat_13804_comb[12]}})) | (p5_bit_slice_13817_comb & {2 {p5_concat_13804_comb[13]}})) | (p5_concat_13818_comb & {2 {p5_concat_13804_comb[14]}})) | (p5_bit_slice_13819_comb & {2 {p5_concat_13804_comb[15]}})) | (p5_bit_slice_13820_comb & {2 {p5_concat_13804_comb[16]}})) | (p5_bit_slice_13821_comb & {2 {p5_concat_13804_comb[17]}})) | (p5_bit_slice_13822_comb & {2 {p5_concat_13804_comb[18]}})) | (p5_bit_slice_13823_comb & {2 {p5_concat_13804_comb[19]}})) | (p5_bit_slice_13824_comb & {2 {p5_concat_13804_comb[20]}})) | (p5_bit_slice_13825_comb & {2 {p5_concat_13804_comb[21]}});
	assign p5_one_hot_sel_14018_comb = ((((((((((((((((((((p5_bit_slice_13827_comb & p5_concat_13826_comb[0]) | (p5_bit_slice_13828_comb & p5_concat_13826_comb[1])) | (p5_bit_slice_13829_comb & p5_concat_13826_comb[2])) | (p5_bit_slice_13830_comb & p5_concat_13826_comb[3])) | (p5_bit_slice_13831_comb & p5_concat_13826_comb[4])) | (p5_bit_slice_13832_comb & p5_concat_13826_comb[5])) | (p5_bit_slice_13737_comb & p5_concat_13826_comb[6])) | (p5_result__10_comb & p5_concat_13826_comb[7])) | (p5_result__39_comb & p5_concat_13826_comb[8])) | (p5_result__32_comb & p5_concat_13826_comb[9])) | (p5_bit_slice_13833_comb & p5_concat_13826_comb[10])) | (p5_bit_slice_13834_comb & p5_concat_13826_comb[11])) | (p5_bit_slice_13835_comb & p5_concat_13826_comb[12])) | (p5_bit_slice_13836_comb & p5_concat_13826_comb[13])) | (p5_bit_slice_13837_comb & p5_concat_13826_comb[14])) | (p5_bit_slice_13838_comb & p5_concat_13826_comb[15])) | (p5_bit_slice_13839_comb & p5_concat_13826_comb[16])) | (p5_bit_slice_13840_comb & p5_concat_13826_comb[17])) | (p5_bit_slice_13841_comb & p5_concat_13826_comb[18])) | (p5_bit_slice_13842_comb & p5_concat_13826_comb[19])) | (p5_bit_slice_13843_comb & p5_concat_13826_comb[20]);
	assign p5_one_hot_sel_14019_comb = (((((((((((((((((((((p5_bit_slice_13844_comb & {6 {p5_concat_13804_comb[0]}}) | (p5_bit_slice_13845_comb & {6 {p5_concat_13804_comb[1]}})) | (p5_bit_slice_13846_comb & {6 {p5_concat_13804_comb[2]}})) | (p5_bit_slice_13847_comb & {6 {p5_concat_13804_comb[3]}})) | (p5_bit_slice_13848_comb & {6 {p5_concat_13804_comb[4]}})) | (p5_bit_slice_13849_comb & {6 {p5_concat_13804_comb[5]}})) | (p5_bit_slice_13850_comb & {6 {p5_concat_13804_comb[6]}})) | (p5_concat_13851_comb & {6 {p5_concat_13804_comb[7]}})) | (p5_bit_slice_13852_comb & {6 {p5_concat_13804_comb[8]}})) | (p5_concat_13853_comb & {6 {p5_concat_13804_comb[9]}})) | (p5_concat_13854_comb & {6 {p5_concat_13804_comb[10]}})) | (p5_bit_slice_13855_comb & {6 {p5_concat_13804_comb[11]}})) | (p5_concat_13856_comb & {6 {p5_concat_13804_comb[12]}})) | (p5_bit_slice_13857_comb & {6 {p5_concat_13804_comb[13]}})) | (p5_bit_slice_13858_comb & {6 {p5_concat_13804_comb[14]}})) | (p5_concat_13859_comb & {6 {p5_concat_13804_comb[15]}})) | (p5_bit_slice_13860_comb & {6 {p5_concat_13804_comb[16]}})) | (p5_bit_slice_13861_comb & {6 {p5_concat_13804_comb[17]}})) | (p5_bit_slice_13862_comb & {6 {p5_concat_13804_comb[18]}})) | (p5_concat_13863_comb & {6 {p5_concat_13804_comb[19]}})) | (p5_bit_slice_13864_comb & {6 {p5_concat_13804_comb[20]}})) | (p5_bit_slice_13865_comb & {6 {p5_concat_13804_comb[21]}});
	assign p5_one_hot_sel_14020_comb = (((((((((((((((((((((p5_bit_slice_13867_comb & {2 {p5_concat_13866_comb[0]}}) | (p5_bit_slice_13868_comb & {2 {p5_concat_13866_comb[1]}})) | (p5_bit_slice_13869_comb & {2 {p5_concat_13866_comb[2]}})) | (p5_bit_slice_13870_comb & {2 {p5_concat_13866_comb[3]}})) | (p5_bit_slice_13871_comb & {2 {p5_concat_13866_comb[4]}})) | (p5_bit_slice_13872_comb & {2 {p5_concat_13866_comb[5]}})) | (p5_concat_13873_comb & {2 {p5_concat_13866_comb[6]}})) | (p5_concat_13874_comb & {2 {p5_concat_13866_comb[7]}})) | (p5_concat_13875_comb & {2 {p5_concat_13866_comb[8]}})) | (p5_concat_13876_comb & {2 {p5_concat_13866_comb[9]}})) | (p5_concat_13877_comb & {2 {p5_concat_13866_comb[10]}})) | (p5_bit_slice_13878_comb & {2 {p5_concat_13866_comb[11]}})) | (p5_bit_slice_13879_comb & {2 {p5_concat_13866_comb[12]}})) | (p5_bit_slice_13880_comb & {2 {p5_concat_13866_comb[13]}})) | (p5_bit_slice_13881_comb & {2 {p5_concat_13866_comb[14]}})) | (p5_bit_slice_13882_comb & {2 {p5_concat_13866_comb[15]}})) | (p5_bit_slice_13883_comb & {2 {p5_concat_13866_comb[16]}})) | (p5_bit_slice_13884_comb & {2 {p5_concat_13866_comb[17]}})) | (p5_bit_slice_13885_comb & {2 {p5_concat_13866_comb[18]}})) | (p5_bit_slice_13886_comb & {2 {p5_concat_13866_comb[19]}})) | (p5_bit_slice_13887_comb & {2 {p5_concat_13866_comb[20]}})) | (p5_bit_slice_13888_comb & {2 {p5_concat_13866_comb[21]}});
	assign p5_one_hot_sel_14021_comb = ((((((((((((((((((((((p5_bit_slice_13890_comb & {2 {p5_concat_13889_comb[0]}}) | (p5_bit_slice_13891_comb & {2 {p5_concat_13889_comb[1]}})) | (p5_bit_slice_13892_comb & {2 {p5_concat_13889_comb[2]}})) | (p5_bit_slice_13893_comb & {2 {p5_concat_13889_comb[3]}})) | (p5_bit_slice_13894_comb & {2 {p5_concat_13889_comb[4]}})) | (p5_bit_slice_13895_comb & {2 {p5_concat_13889_comb[5]}})) | (p5_bit_slice_13896_comb & {2 {p5_concat_13889_comb[6]}})) | (p5_bit_slice_13897_comb & {2 {p5_concat_13889_comb[7]}})) | (p5_concat_13898_comb & {2 {p5_concat_13889_comb[8]}})) | (p5_bit_slice_13899_comb & {2 {p5_concat_13889_comb[9]}})) | (p5_concat_13900_comb & {2 {p5_concat_13889_comb[10]}})) | (p5_concat_13901_comb & {2 {p5_concat_13889_comb[11]}})) | (p5_bit_slice_13902_comb & {2 {p5_concat_13889_comb[12]}})) | (p5_bit_slice_13903_comb & {2 {p5_concat_13889_comb[13]}})) | (p5_bit_slice_13904_comb & {2 {p5_concat_13889_comb[14]}})) | (p5_concat_13905_comb & {2 {p5_concat_13889_comb[15]}})) | (p5_bit_slice_13906_comb & {2 {p5_concat_13889_comb[16]}})) | (p5_bit_slice_13907_comb & {2 {p5_concat_13889_comb[17]}})) | (p5_bit_slice_13908_comb & {2 {p5_concat_13889_comb[18]}})) | (p5_bit_slice_13909_comb & {2 {p5_concat_13889_comb[19]}})) | (p5_xor_13910_comb & {2 {p5_concat_13889_comb[20]}})) | (p5_bit_slice_13911_comb & {2 {p5_concat_13889_comb[21]}})) | (p5_bit_slice_13912_comb & {2 {p5_concat_13889_comb[22]}});
	assign p5_one_hot_sel_14022_comb = (((((((((((((((((((((p5_bit_slice_13914_comb & {4 {p5_concat_13913_comb[0]}}) | (p5_bit_slice_13915_comb & {4 {p5_concat_13913_comb[1]}})) | (p5_bit_slice_13916_comb & {4 {p5_concat_13913_comb[2]}})) | (p5_bit_slice_13917_comb & {4 {p5_concat_13913_comb[3]}})) | (p5_bit_slice_13918_comb & {4 {p5_concat_13913_comb[4]}})) | (p5_bit_slice_13919_comb & {4 {p5_concat_13913_comb[5]}})) | (p5_bit_slice_13920_comb & {4 {p5_concat_13913_comb[6]}})) | (p5_bit_slice_13921_comb & {4 {p5_concat_13913_comb[7]}})) | (p5_concat_13922_comb & {4 {p5_concat_13913_comb[8]}})) | (p5_bit_slice_13923_comb & {4 {p5_concat_13913_comb[9]}})) | (p5_concat_13924_comb & {4 {p5_concat_13913_comb[10]}})) | (p5_concat_13925_comb & {4 {p5_concat_13913_comb[11]}})) | (p5_bit_slice_13926_comb & {4 {p5_concat_13913_comb[12]}})) | (p5_concat_13927_comb & {4 {p5_concat_13913_comb[13]}})) | (p5_bit_slice_13928_comb & {4 {p5_concat_13913_comb[14]}})) | (p5_bit_slice_13929_comb & {4 {p5_concat_13913_comb[15]}})) | (p5_bit_slice_13930_comb & {4 {p5_concat_13913_comb[16]}})) | (p5_bit_slice_13931_comb & {4 {p5_concat_13913_comb[17]}})) | (p5_bit_slice_13932_comb & {4 {p5_concat_13913_comb[18]}})) | (p5_bit_slice_13933_comb & {4 {p5_concat_13913_comb[19]}})) | (p5_bit_slice_13934_comb & {4 {p5_concat_13913_comb[20]}})) | (p5_bit_slice_13935_comb & {4 {p5_concat_13913_comb[21]}});
	assign p5_one_hot_sel_14023_comb = ((((((((((((((((((((p5_bit_slice_13937_comb & p5_concat_13936_comb[0]) | (p5_bit_slice_13938_comb & p5_concat_13936_comb[1])) | (p5_bit_slice_13939_comb & p5_concat_13936_comb[2])) | (p5_bit_slice_13940_comb & p5_concat_13936_comb[3])) | (p5_bit_slice_13941_comb & p5_concat_13936_comb[4])) | (p5_bit_slice_13942_comb & p5_concat_13936_comb[5])) | (p5_result__25_comb & p5_concat_13936_comb[6])) | (p5_bit_slice_13735_comb & p5_concat_13936_comb[7])) | (p5_result__39_comb & p5_concat_13936_comb[8])) | (p5_result__10_comb & p5_concat_13936_comb[9])) | (p5_result__17_comb & p5_concat_13936_comb[10])) | (p5_bit_slice_13943_comb & p5_concat_13936_comb[11])) | (p5_bit_slice_13944_comb & p5_concat_13936_comb[12])) | (p5_bit_slice_13945_comb & p5_concat_13936_comb[13])) | (p5_bit_slice_13946_comb & p5_concat_13936_comb[14])) | (p5_bit_slice_13947_comb & p5_concat_13936_comb[15])) | (p5_bit_slice_13948_comb & p5_concat_13936_comb[16])) | (p5_bit_slice_13949_comb & p5_concat_13936_comb[17])) | (p5_bit_slice_13950_comb & p5_concat_13936_comb[18])) | (p5_bit_slice_13951_comb & p5_concat_13936_comb[19])) | (p5_bit_slice_13952_comb & p5_concat_13936_comb[20]);
	assign p5_one_hot_sel_14024_comb = ((((((((((((((((((((p5_bit_slice_13954_comb & {5 {p5_concat_13953_comb[0]}}) | (p5_bit_slice_13955_comb & {5 {p5_concat_13953_comb[1]}})) | (p5_bit_slice_13956_comb & {5 {p5_concat_13953_comb[2]}})) | (p5_bit_slice_13957_comb & {5 {p5_concat_13953_comb[3]}})) | (p5_bit_slice_13958_comb & {5 {p5_concat_13953_comb[4]}})) | (p5_bit_slice_13959_comb & {5 {p5_concat_13953_comb[5]}})) | (p5_bit_slice_13960_comb & {5 {p5_concat_13953_comb[6]}})) | (p5_concat_13961_comb & {5 {p5_concat_13953_comb[7]}})) | (p5_bit_slice_13594_comb & {5 {p5_concat_13953_comb[8]}})) | (p5_concat_13962_comb & {5 {p5_concat_13953_comb[9]}})) | (p5_concat_13963_comb & {5 {p5_concat_13953_comb[10]}})) | (p5_concat_13964_comb & {5 {p5_concat_13953_comb[11]}})) | (p5_bit_slice_13965_comb & {5 {p5_concat_13953_comb[12]}})) | (p5_bit_slice_13966_comb & {5 {p5_concat_13953_comb[13]}})) | (p5_bit_slice_13967_comb & {5 {p5_concat_13953_comb[14]}})) | (p5_concat_13968_comb & {5 {p5_concat_13953_comb[15]}})) | (p5_bit_slice_13969_comb & {5 {p5_concat_13953_comb[16]}})) | (p5_bit_slice_13970_comb & {5 {p5_concat_13953_comb[17]}})) | (p5_bit_slice_13971_comb & {5 {p5_concat_13953_comb[18]}})) | (p5_bit_slice_13972_comb & {5 {p5_concat_13953_comb[19]}})) | (p5_bit_slice_13973_comb & {5 {p5_concat_13953_comb[20]}});
	assign p5_one_hot_sel_14025_comb = (((((((((((((((((((((p5_bit_slice_13975_comb & {2 {p5_concat_13974_comb[0]}}) | (p5_bit_slice_13976_comb & {2 {p5_concat_13974_comb[1]}})) | (p5_bit_slice_13977_comb & {2 {p5_concat_13974_comb[2]}})) | (p5_bit_slice_13978_comb & {2 {p5_concat_13974_comb[3]}})) | (p5_bit_slice_13979_comb & {2 {p5_concat_13974_comb[4]}})) | (p5_bit_slice_13980_comb & {2 {p5_concat_13974_comb[5]}})) | (p5_bit_slice_13981_comb & {2 {p5_concat_13974_comb[6]}})) | (p5_concat_13982_comb & {2 {p5_concat_13974_comb[7]}})) | (p5_bit_slice_13983_comb & {2 {p5_concat_13974_comb[8]}})) | (p5_concat_13984_comb & {2 {p5_concat_13974_comb[9]}})) | (p5_concat_13985_comb & {2 {p5_concat_13974_comb[10]}})) | (p5_bit_slice_13986_comb & {2 {p5_concat_13974_comb[11]}})) | (p5_bit_slice_13987_comb & {2 {p5_concat_13974_comb[12]}})) | (p5_bit_slice_13988_comb & {2 {p5_concat_13974_comb[13]}})) | (p5_bit_slice_13989_comb & {2 {p5_concat_13974_comb[14]}})) | (p5_bit_slice_13990_comb & {2 {p5_concat_13974_comb[15]}})) | (p5_bit_slice_13991_comb & {2 {p5_concat_13974_comb[16]}})) | (p5_bit_slice_13992_comb & {2 {p5_concat_13974_comb[17]}})) | (p5_bit_slice_13993_comb & {2 {p5_concat_13974_comb[18]}})) | (p5_bit_slice_13994_comb & {2 {p5_concat_13974_comb[19]}})) | (p5_bit_slice_13995_comb & {2 {p5_concat_13974_comb[20]}})) | (p5_bit_slice_13996_comb & {2 {p5_concat_13974_comb[21]}});
	assign p5_one_hot_sel_14026_comb = (((((((((((((((((((p5_bit_slice_13998_comb & p5_concat_13997_comb[0]) | (p5_bit_slice_13999_comb & p5_concat_13997_comb[1])) | (p5_bit_slice_14000_comb & p5_concat_13997_comb[2])) | (p5_bit_slice_14001_comb & p5_concat_13997_comb[3])) | (p5_bit_slice_14002_comb & p5_concat_13997_comb[4])) | (p5_bit_slice_14003_comb & p5_concat_13997_comb[5])) | (p5_rotation_1__6_comb & p5_concat_13997_comb[6])) | (p5_result__23_comb & p5_concat_13997_comb[7])) | (p5_result__26_comb & p5_concat_13997_comb[8])) | (p5_bit_slice_14004_comb & p5_concat_13997_comb[9])) | (p5_bit_slice_14005_comb & p5_concat_13997_comb[10])) | (p5_bit_slice_14006_comb & p5_concat_13997_comb[11])) | (p5_bit_slice_14007_comb & p5_concat_13997_comb[12])) | (p5_bit_slice_14008_comb & p5_concat_13997_comb[13])) | (p5_bit_slice_14009_comb & p5_concat_13997_comb[14])) | (p5_bit_slice_14010_comb & p5_concat_13997_comb[15])) | (p5_bit_slice_14011_comb & p5_concat_13997_comb[16])) | (p5_bit_slice_14012_comb & p5_concat_13997_comb[17])) | (p5_bit_slice_14013_comb & p5_concat_13997_comb[18])) | (p5_bit_slice_14014_comb & p5_concat_13997_comb[19]);
	assign p5_concat_14027_comb = {p5_one_hot_sel_14015_comb, p5_one_hot_sel_14016_comb, p5_one_hot_sel_14017_comb, p5_one_hot_sel_14018_comb, p5_one_hot_sel_14019_comb, p5_one_hot_sel_14020_comb, p5_one_hot_sel_14021_comb, p5_one_hot_sel_14022_comb, p5_one_hot_sel_14023_comb, p5_one_hot_sel_14024_comb, p5_one_hot_sel_14025_comb, p5_one_hot_sel_14026_comb};
	assign p5_sign_ext_14028_comb = {32 {p4_valid}};
	assign p5_and_14029_comb = p5_concat_14027_comb & p5_sign_ext_14028_comb;
	assign p5_tuple_14030_comb = {p4_and_13245, p5_and_14029_comb};
	reg [32:0] p5_tuple_14030;
	always @(posedge clk) p5_tuple_14030 <= p5_tuple_14030_comb;
	assign out = p5_tuple_14030;
endmodule
